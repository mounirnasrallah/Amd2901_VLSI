* Spice description of amd2901
* Spice driver version 1074415736
* Date ( dd/mm/yyyy hh:mm:ss ): 10/06/2014 at  1:31:03

* INTERF a[0] a[1] a[2] a[3] b[0] b[1] b[2] b[3] cin clk cout d[0] d[1] d[2] 
* INTERF d[3] f3 i[0] i[1] i[2] i[3] i[4] i[5] i[6] i[7] i[8] ng noe np ovr 
* INTERF q0 q3 r0 r3 vdde vddi vsse vssi y[0] y[1] y[2] y[3] zero 


.subckt amd2901 3662 3136 2467 1941 1402 735 177 159 4408 180 4400 4545 4544 
+ 4543 4542 151 44 39 34 29 24 19 14 9 4 3573 738 3027 1828 4125 4128 4380 
+ 4371 4535 4478 4541 4540 4539 4538 4537 4536 1280 
* NET 1 = p_i8.node_cp
* NET 3 = p_i8.n6d
* NET 4 = i[8]
* NET 5 = p_i8.1019ymous_
* NET 6 = p_i7.585nymous_
* NET 7 = p_i7.31onymous_
* NET 8 = p_i7.n6d
* NET 9 = i[7]
* NET 10 = p_i7.vdde
* NET 11 = p_i6.node_cp
* NET 13 = p_i6.n6d
* NET 14 = i[6]
* NET 15 = p_i6.903nymous_
* NET 16 = p_i5.node_cp
* NET 18 = p_i5.n6d
* NET 19 = i[5]
* NET 20 = p_i5.1019ymous_
* NET 21 = p_i4.node_cp
* NET 23 = p_i4.n6d
* NET 24 = i[4]
* NET 25 = p_i4.1019ymous_
* NET 26 = p_i3.585nymous_
* NET 27 = p_i3.405nymous_
* NET 28 = p_i3.n6d
* NET 29 = i[3]
* NET 30 = p_i3.vdde
* NET 31 = p_i2.node_cp
* NET 33 = p_i2.312nymous_
* NET 34 = i[2]
* NET 35 = p_i2.903nymous_
* NET 36 = p_i1.node_cp
* NET 38 = p_i1.312nymous_
* NET 39 = i[1]
* NET 40 = p_i1.1019ymous_
* NET 41 = p_i0.585nymous_
* NET 43 = p_i0.n6d
* NET 44 = i[0]
* NET 45 = p_i0.vdde
* NET 46 = p_i8.766nymous_
* NET 47 = p_i8.n1
* NET 48 = p_i8.n0
* NET 49 = p_i8.79onymous_
* NET 50 = p_i8.58onymous_
* NET 51 = p_i8.n16c
* NET 52 = p_i8.nnt
* NET 53 = p_i8.1066ymous_
* NET 54 = p_i7.n5b
* NET 55 = p_i7.n0
* NET 56 = p_i7.79onymous_
* NET 57 = p_i7.93onymous_
* NET 58 = p_i7.58onymous_
* NET 59 = p_i7.n16c
* NET 60 = p_i7.259nymous_
* NET 61 = p_i7.196nymous_
* NET 62 = p_i6.n5a
* NET 63 = p_i6.111nymous_
* NET 64 = p_i6.n1
* NET 65 = p_i6.42onymous_
* NET 66 = p_i6.58onymous_
* NET 67 = p_i6.n16a
* NET 68 = p_i6.nnt
* NET 69 = p_i6.nt
* NET 70 = p_i5.766nymous_
* NET 71 = p_i5.n1
* NET 72 = p_i5.n0
* NET 73 = p_i5.79onymous_
* NET 74 = p_i5.58onymous_
* NET 75 = p_i5.n16c
* NET 76 = p_i5.259nymous_
* NET 77 = p_i5.1066ymous_
* NET 78 = p_vddeck1.246nymous_
* NET 79 = p_vddeck1.64onymous_
* NET 80 = p_vddeck0.253nymous_
* NET 81 = p_vddeck0.64onymous_
* NET 82 = p_i4.766nymous_
* NET 83 = p_i4.n1
* NET 84 = p_i4.n0
* NET 85 = p_i4.79onymous_
* NET 86 = p_i4.58onymous_
* NET 87 = p_i4.n16c
* NET 88 = p_i4.259nymous_
* NET 89 = p_i4.1066ymous_
* NET 90 = p_i3.n5b
* NET 91 = p_i3.n0
* NET 92 = p_i3.n4b
* NET 93 = p_i3.79onymous_
* NET 94 = p_i3.93onymous_
* NET 95 = p_i3.n16c
* NET 96 = p_i3.259nymous_
* NET 97 = p_i3.196nymous_
* NET 98 = p_i2.n5a
* NET 99 = p_i2.111nymous_
* NET 100 = p_i2.n1
* NET 101 = p_i2.42onymous_
* NET 102 = p_i2.58onymous_
* NET 103 = p_i2.n16a
* NET 104 = p_i2.nnt
* NET 105 = p_i2.nt
* NET 106 = p_i1.766nymous_
* NET 107 = p_i1.n1
* NET 108 = p_i1.n0
* NET 109 = p_i1.532nymous_
* NET 111 = p_i1.n16a
* NET 112 = p_i1.259nymous_
* NET 113 = p_i1.1066ymous_
* NET 114 = p_i0.160nymous_
* NET 115 = p_i0.n0
* NET 116 = p_i0.79onymous_
* NET 117 = p_i0.58onymous_
* NET 118 = p_i0.n1
* NET 119 = p_i0.n16c
* NET 120 = p_i0.259nymous_
* NET 121 = p_i0.221nymous_
* NET 122 = p_i8.1061ymous_
* NET 123 = i_from_pads[7]
* NET 124 = p_i6.1061ymous_
* NET 125 = p_i5.1060ymous_
* NET 126 = p_vddeck1.cko
* NET 127 = p_vddeck0.cko
* NET 128 = p_i4.1060ymous_
* NET 130 = i_from_pads[3]
* NET 131 = p_i0.1060ymous_
* NET 132 = p_f3.137nymous_
* NET 133 = p_b3.639nymous_
* NET 134 = p_b3.132nymous_
* NET 135 = p_f3.69onymous_
* NET 136 = p_f3.n17a
* NET 137 = p_b3.p1
* NET 138 = p_b3.57onymous_
* NET 139 = p_f3.n16b
* NET 140 = p_b3.1280ymous_
* NET 141 = p_b3.cpb
* NET 142 = p_b3.324nymous_
* NET 144 = p_f3.p6c
* NET 145 = p_f3.301nymous_
* NET 146 = p_f3.305nymous_
* NET 147 = p_f3.274nymous_
* NET 148 = f3_to_pads
* NET 149 = p_b3.nnt
* NET 150 = p_f3.227nymous_
* NET 151 = f3
* NET 152 = p_f3.197nymous_
* NET 153 = p_f3.224nymous_
* NET 154 = p_f3.193nymous_
* NET 155 = p_b3.1066ymous_
* NET 156 = p_b3.197nymous_
* NET 157 = p_b3.n14c
* NET 159 = b[3]
* NET 160 = p_f3.318nymous_
* NET 161 = p_b2.132nymous_
* NET 162 = p_b2.93onymous_
* NET 163 = p_b2.p2
* NET 164 = p_b2.cpb
* NET 165 = p_b2.414nymous_
* NET 166 = p_b2.n8b
* NET 168 = p_ck.p6a
* NET 169 = p_ck.24onymous_
* NET 170 = p_b2.259nymous_
* NET 171 = p_b2.1280ymous_
* NET 172 = p_ck.507nymous_
* NET 173 = p_ck.115nymous_
* NET 175 = p_b2.196nymous_
* NET 176 = b_from_pads[2]
* NET 177 = b[2]
* NET 178 = p_ck.711nymous_
* NET 179 = p_ck.720nymous_
* NET 180 = clk
* NET 200 = p_b2.n14a
* NET 201 = p_b2.568nymous_
* NET 207 = core.iram.not_aux144
* NET 210 = core.iram.not_aux144_ins.i0
* NET 211 = core.iram.inv_x2_3_sig
* NET 212 = core.iram.aux99_ins.i1
* NET 213 = b_from_pads[0]
* NET 229 = core.iram.not_aux84
* NET 238 = core.iram.not_aux52
* NET 245 = core.iram.ab_data_idx_10_1_ins.sff_m
* NET 247 = core.iram.ab_data_idx_10_1_ins.y
* NET 248 = core.iram.ab_data_idx_10_1_ins.sff_s
* NET 249 = core.iram.ab_data_idx_10_1_ins.ck
* NET 250 = core.iram.ab_data_idx_10_1_ins.nckr
* NET 251 = core.iram.ab_data_idx_10_1_ins.u
* NET 253 = core.iram.ab_data_idx_10_1_ins.ckr
* NET 255 = core.iram.na2_x1_40_sig
* NET 258 = core.iram.ao22_x2_38_sig
* NET 265 = core.iram.not_aux31
* NET 271 = core.iram.ab_data_idx_1_2_ins.sff_s
* NET 272 = core.iram.ab_data_idx_1_2_ins.y
* NET 274 = core.iram.ab_data_idx_1_2_ins.u
* NET 275 = core.iram.ab_data_idx_1_2_ins.sff_m
* NET 278 = core.iram.ab_data_idx_1_2_ins.nckr
* NET 280 = core.iram.ab_data_idx_1_2_ins.ckr
* NET 283 = core.iram.ao22_x2_7_sig
* NET 288 = core.iram.na2_x1_9_sig
* NET 291 = core.iram.not_aux53
* NET 296 = core.iram.not_aux54
* NET 300 = core.iram.not_aux33_ins.i0
* NET 303 = core.iram.not_aux32
* NET 309 = core.iram.ab_data_idx_0_2_ins.y
* NET 310 = core.iram.ab_data_idx_0_2_ins.sff_s
* NET 312 = core.iram.ab_data_idx_0_2_ins.sff_m
* NET 314 = core.iram.ab_data_idx_0_2_ins.ck
* NET 315 = core.iram.ab_data_idx_0_2_ins.u
* NET 317 = core.iram.ab_data_idx_0_2_ins.ckr
* NET 320 = core.iram.ao22_x2_3_sig
* NET 321 = core.iram.ab_data_idx_0_2_ins.nckr
* NET 326 = core.iram.na2_x1_5_sig
* NET 328 = core.iram.not_aux33
* NET 332 = core.iram.not_aux64
* NET 335 = core.iram.na2_x1_17_sig
* NET 341 = core.iram.ab_data_idx_3_2_ins.sff_s
* NET 342 = core.iram.ao22_x2_15_sig
* NET 343 = core.iram.ab_data_idx_3_2_ins.y
* NET 348 = core.iram.ab_data_idx_3_2_ins.sff_m
* NET 350 = core.iram.ab_data_idx_3_2_ins.ckr
* NET 351 = core.iram.ab_data_idx_3_2_ins.nckr
* NET 352 = core.iram.ab_data_idx_3_2_ins.u
* NET 353 = core.iram.ab_data_idx_15_1_ins.sff_s
* NET 356 = core.iram.ab_data_idx_15_1_ins.y
* NET 358 = core.iram.ab_data_idx_15_1_ins.sff_m
* NET 359 = core.iram.ab_data_idx_15_1_ins.ck
* NET 360 = core.iram.ab_data_idx_15_1_ins.nckr
* NET 361 = core.iram.ab_data_idx_15_1_ins.u
* NET 362 = core.iram.ab_data_idx_15_1_ins.ckr
* NET 363 = core.iram.aux97_ins.i0
* NET 365 = core.iram.aux97
* NET 367 = core.iram.not_b_0_ins.i
* NET 369 = core.iram.ab_data_idx_9_2_ins.sff_s
* NET 370 = core.iram.ab_data_idx_9_2_ins.y
* NET 372 = core.iram.ab_data_idx_9_2_ins.u
* NET 374 = core.iram.ab_data_idx_9_2_ins.sff_m
* NET 375 = core.iram.a3_x2_3_sig
* NET 377 = core.iram.ab_data_idx_9_2_ins.ckr
* NET 378 = core.iram.ab_data_idx_9_2_ins.nckr
* NET 380 = core.iram.noa22_x1_2_sig
* NET 381 = core.iram.inv_x2_6_sig
* NET 385 = core.iram.not_aux74
* NET 388 = core.iram.ab_data_idx_8_2_ins.sff_s
* NET 389 = core.iram.ab_data_idx_8_2_ins.y
* NET 391 = core.iram.ab_data_idx_8_2_ins.sff_m
* NET 392 = core.iram.ab_data_idx_8_2_ins.ck
* NET 393 = core.iram.ab_data_idx_8_2_ins.u
* NET 395 = core.iram.ab_data_idx_8_2_ins.ckr
* NET 396 = core.iram.ab_data_idx_8_2_ins.nckr
* NET 397 = core.iram.ao22_x2_35_sig
* NET 400 = core.iram.na2_x1_37_sig
* NET 402 = core.iram.not_aux77
* NET 404 = core.iram.not_aux76
* NET 406 = core.iram.not_aux22
* NET 409 = core.iram.na2_x1_41_sig
* NET 412 = core.iram.ab_data_idx_10_2_ins.y
* NET 415 = core.iram.ab_data_idx_10_2_ins.sff_s
* NET 416 = core.iram.ao22_x2_39_sig
* NET 417 = core.iram.ab_data_idx_10_2_ins.ckr
* NET 418 = core.iram.ab_data_idx_10_2_ins.u
* NET 420 = core.iram.ab_data_idx_10_2_ins.sff_m
* NET 422 = core.iram.ab_data_idx_10_2_ins.nckr
* NET 424 = core.iram.ab_data_idx_0_1_ins.sff_s
* NET 426 = core.iram.ab_data_idx_0_1_ins.y
* NET 428 = core.iram.ab_data_idx_0_1_ins.sff_m
* NET 429 = core.iram.ab_data_idx_0_1_ins.u
* NET 431 = p_noe.1061ymous_
* NET 432 = core.iram.ab_data_idx_0_1_ins.ck
* NET 433 = core.iram.ab_data_idx_0_1_ins.nckr
* NET 434 = core.iram.ab_data_idx_0_1_ins.ckr
* NET 435 = core.iram.ao22_x2_2_sig
* NET 438 = core.iram.not_aux24_ins.i0
* NET 440 = core.iram.na2_x1_4_sig
* NET 441 = core.iram.not_aux24
* NET 444 = core.iram.ab_data_idx_3_1_ins.sff_s
* NET 445 = core.iram.ab_data_idx_3_1_ins.y
* NET 447 = core.iram.ab_data_idx_3_1_ins.sff_m
* NET 449 = core.iram.ab_data_idx_3_1_ins.nckr
* NET 450 = core.iram.ab_data_idx_3_1_ins.u
* NET 451 = core.iram.ab_data_idx_3_1_ins.ckr
* NET 452 = core.iram.na2_x1_16_sig
* NET 455 = core.iram.ao22_x2_14_sig
* NET 458 = core.iram.na2_x1_33_sig
* NET 463 = core.iram.ab_data_idx_7_2_ins.sff_s
* NET 464 = core.iram.ao22_x2_31_sig
* NET 465 = core.iram.ab_data_idx_7_2_ins.y
* NET 468 = core.iram.ab_data_idx_7_2_ins.sff_m
* NET 469 = core.iram.ab_data_idx_7_2_ins.ck
* NET 470 = core.iram.ab_data_idx_7_2_ins.u
* NET 471 = core.iram.ab_data_idx_7_2_ins.nckr
* NET 472 = core.iram.ab_data_idx_7_2_ins.ckr
* NET 473 = p_b1.112nymous_
* NET 474 = p_b1.640nymous_
* NET 475 = p_noe.n17d
* NET 479 = core.iram.aux99_ins.nq
* NET 506 = p_b1.43onymous_
* NET 507 = p_b1.466nymous_
* NET 508 = p_noe.25onymous_
* NET 510 = core.iram.a2_x2_3_sig
* NET 511 = core.iram.oa2ao222_x2_2_sig
* NET 515 = core.iram.nao22_x1_7_ins.i0
* NET 516 = core.iram.nao22_x1_7_sig
* NET 520 = core.iram.not_b_3_ins.i
* NET 521 = core.iram.not_ab_data_idx_15[1]
* NET 527 = core.iram.ab_data_idx_8_1_ins.sff_m
* NET 528 = core.iram.ab_data_idx_8_1_ins.y
* NET 529 = core.iram.ab_data_idx_8_1_ins.sff_s
* NET 533 = core.iram.ab_data_idx_8_1_ins.u
* NET 535 = core.iram.ab_data_idx_8_1_ins.ckr
* NET 536 = core.iram.ab_data_idx_8_1_ins.nckr
* NET 537 = core.iram.not_aux134
* NET 544 = core.iram.not_aux83
* NET 547 = core.iram.ao22_x2_34_sig
* NET 553 = core.iram.na2_x1_36_sig
* NET 555 = core.iram.not_aux75
* NET 561 = core.iram.ab_data_idx_12_2_ins.sff_m
* NET 563 = core.iram.ab_data_idx_12_2_ins.y
* NET 564 = core.iram.ab_data_idx_12_2_ins.sff_s
* NET 566 = core.iram.ab_data_idx_12_2_ins.ck
* NET 567 = core.iram.ab_data_idx_12_2_ins.nckr
* NET 568 = core.iram.ab_data_idx_12_2_ins.u
* NET 569 = core.iram.ab_data_idx_12_2_ins.ckr
* NET 572 = core.iram.na2_x1_45_sig
* NET 573 = core.iram.ao22_x2_43_sig
* NET 576 = core.iram.not_aux88
* NET 581 = core.iram.not_aux49
* NET 589 = core.iram.ab_data_idx_1_1_ins.sff_s
* NET 591 = core.iram.ab_data_idx_1_1_ins.sff_m
* NET 593 = core.iram.ab_data_idx_1_1_ins.y
* NET 597 = core.iram.ab_data_idx_1_1_ins.u
* NET 598 = core.iram.ab_data_idx_1_1_ins.ckr
* NET 599 = core.iram.ab_data_idx_1_1_ins.nckr
* NET 600 = core.iram.ao22_x2_6_sig
* NET 603 = core.iram.na2_x1_8_sig
* NET 605 = core.iram.not_aux50
* NET 608 = core.iram.not_aux51_ins.i0
* NET 614 = core.iram.not_aux51
* NET 616 = core.iram.ab_data_idx_5_1_ins.y
* NET 617 = core.iram.ab_data_idx_5_1_ins.sff_s
* NET 620 = core.iram.ab_data_idx_5_1_ins.u
* NET 622 = core.iram.ab_data_idx_5_1_ins.sff_m
* NET 624 = core.iram.ab_data_idx_5_1_ins.ckr
* NET 625 = core.iram.ab_data_idx_5_1_ins.ck
* NET 626 = core.iram.ao22_x2_22_sig
* NET 627 = core.iram.ab_data_idx_5_1_ins.nckr
* NET 630 = core.iram.na2_x1_24_sig
* NET 633 = core.iram.not_aux23
* NET 637 = core.iram.ab_data_idx_4_1_ins.sff_s
* NET 640 = core.iram.ab_data_idx_4_1_ins.y
* NET 641 = core.iram.ab_data_idx_4_1_ins.sff_m
* NET 646 = core.iram.ab_data_idx_4_1_ins.ckr
* NET 647 = core.iram.ab_data_idx_4_1_ins.nckr
* NET 648 = core.iram.ab_data_idx_4_1_ins.u
* NET 649 = core.iram.na2_x1_20_sig
* NET 651 = core.iram.ao22_x2_18_sig
* NET 654 = core.iram.na2_x1_21_sig
* NET 658 = core.iram.not_aux63
* NET 661 = core.iram.not_aux59
* NET 662 = core.iram.na2_x1_32_sig
* NET 667 = core.iram.ab_data_idx_7_1_ins.sff_s
* NET 669 = core.iram.ao22_x2_30_sig
* NET 670 = core.iram.ab_data_idx_7_1_ins.y
* NET 673 = core.iram.ab_data_idx_7_1_ins.sff_m
* NET 676 = core.iram.ab_data_idx_7_1_ins.ck
* NET 677 = core.iram.ab_data_idx_7_1_ins.ckr
* NET 678 = core.iram.ab_data_idx_7_1_ins.nckr
* NET 679 = core.iram.ab_data_idx_7_1_ins.u
* NET 680 = p_b1.n6a
* NET 681 = p_b1.1280ymous_
* NET 682 = p_b1.n8a
* NET 683 = p_b1.324nymous_
* NET 684 = p_noe.p6a
* NET 686 = p_noe.p7a
* NET 687 = p_noe.n2
* NET 688 = p_noe.129nymous_
* NET 689 = core.iram.a2_x2_4_ins.i1
* NET 692 = core.iram.na3_x1_5_sig
* NET 693 = core.iram.not_aux145
* NET 694 = core.iram.na3_x1_6_sig
* NET 696 = core.iram.inv_x2_9_sig
* NET 700 = core.iram.ab_data_idx_12_1_ins.ck
* NET 701 = core.iram.na2_x1_44_sig
* NET 703 = core.iram.not_aux11_ins.i0
* NET 704 = core.iram.not_aux11_ins.i1
* NET 706 = core.iram.aux109
* NET 707 = a_from_pads[1]
* NET 708 = core.iram.ab_data_idx_9[2]
* NET 709 = core.iram.na3_x1_23_sig
* NET 710 = core.iram.na3_x1_24_sig
* NET 713 = core.iram.na3_x1_25_sig
* NET 714 = core.iram.na3_x1_24_ins.i0
* NET 715 = core.iram.ab_data_idx_1[2]
* NET 716 = core.iram.na3_x1_58_sig
* NET 720 = core.iram.na3_x1_57_ins.i0
* NET 721 = core.iram.na3_x1_57_sig
* NET 723 = core.iram.ab_data_idx_0[2]
* NET 725 = core.iram.na3_x1_55_sig
* NET 728 = core.iram.not_aux58
* NET 730 = core.iram.ao22_x2_31_ins.i1
* NET 731 = core.iram.aux62_ins.i0
* NET 733 = core.iram.ab_data_idx_6_2_ins.ck
* NET 734 = p_b1.nnt
* NET 735 = b[1]
* NET 736 = p_noe.772nymous_
* NET 737 = p_noe.815nymous_
* NET 738 = noe
* NET 739 = p_noe.156nymous_
* NET 740 = p_noe.766nymous_
* NET 743 = core.iram.a2_x2_4_sig
* NET 745 = core.iram.a2_x2_2_sig
* NET 748 = core.iram.ab_data_idx_11_1_ins.ckr
* NET 749 = core.iram.ab_data_idx_11_1_ins.nckr
* NET 750 = core.iram.ab_data_idx_11_1_ins.sff_m
* NET 751 = core.iram.ab_data_idx_11_1_ins.y
* NET 753 = core.iram.ab_data_idx_11_1_ins.sff_s
* NET 755 = core.iram.noa2a22_x1_3_sig
* NET 758 = core.iram.ab_data_idx_11_1_ins.u
* NET 763 = core.iram.not_aux117
* NET 765 = core.iram.not_aux125
* NET 766 = core.iram.ab_data_idx_12_1_ins.ckr
* NET 767 = core.iram.ab_data_idx_12_1_ins.nckr
* NET 768 = core.iram.ab_data_idx_12_1_ins.sff_m
* NET 769 = core.iram.ab_data_idx_12_1_ins.y
* NET 771 = core.iram.ab_data_idx_12_1_ins.sff_s
* NET 774 = core.iram.ab_data_idx_12_1_ins.u
* NET 777 = core.iram.ao22_x2_42_sig
* NET 785 = core.iram.not_aux11
* NET 787 = core.iram.ab_data_idx_4_2_ins.ckr
* NET 788 = core.iram.ab_data_idx_4_2_ins.nckr
* NET 791 = core.iram.ab_data_idx_4_2_ins.sff_s
* NET 792 = core.iram.ab_data_idx_4_2_ins.sff_m
* NET 794 = core.iram.ab_data_idx_4_2_ins.y
* NET 796 = core.iram.ao22_x2_19_sig
* NET 799 = core.iram.ab_data_idx_4_2_ins.u
* NET 803 = core.iram.aux157
* NET 807 = core.iram.ab_data_idx_6_2_ins.ckr
* NET 808 = core.iram.ab_data_idx_6_2_ins.nckr
* NET 809 = core.iram.ab_data_idx_6_2_ins.sff_s
* NET 812 = core.iram.ab_data_idx_6_2_ins.y
* NET 813 = core.iram.ab_data_idx_6_2_ins.sff_m
* NET 818 = core.iram.ab_data_idx_6_2_ins.u
* NET 819 = p_b1.nt
* NET 820 = p_b1.970nymous_
* NET 821 = p_b1.n14b
* NET 822 = p_b1.87onymous_
* NET 825 = core.iram.inv_x2_sig
* NET 829 = core.iram.aux139
* NET 830 = core.iram.na4_x1_ins.i2
* NET 835 = core.iram.ab_data_idx_9_1_ins.y
* NET 836 = core.iram.ab_data_idx_9_1_ins.sff_s
* NET 837 = core.iram.ab_data_idx_9_1_ins.sff_m
* NET 840 = core.iram.ab_data_idx_9_1_ins.u
* NET 842 = core.iram.ab_data_idx_9_1_ins.ckr
* NET 843 = core.iram.a3_x2_2_sig
* NET 844 = core.iram.ab_data_idx_9_1_ins.nckr
* NET 845 = core.iram.noa22_x1_sig
* NET 846 = core.iram.inv_x2_5_sig
* NET 848 = core.iram.not_aux118_ins.i0
* NET 853 = core.iram.not_aux126
* NET 855 = core.iram.not_aux118
* NET 856 = core.iram.not_aux92
* NET 859 = core.iram.inv_x2_10_sig
* NET 861 = core.iram.ab_data_idx_11_2_ins.sff_s
* NET 862 = core.iram.ab_data_idx_11_2_ins.y
* NET 864 = core.iram.ab_data_idx_11_2_ins.sff_m
* NET 866 = core.iram.ab_data_idx_11_2_ins.ck
* NET 867 = core.iram.noa2a22_x1_4_sig
* NET 868 = core.iram.ab_data_idx_11_2_ins.u
* NET 869 = core.iram.ab_data_idx_11_2_ins.ckr
* NET 870 = core.iram.ab_data_idx_11_2_ins.nckr
* NET 871 = core.iram.na3_x1_47_sig
* NET 874 = core.iram.na3_x1_46_sig
* NET 877 = core.iram.ab_data_idx_9[1]
* NET 882 = core.iram.na3_x1_56_sig
* NET 884 = core.iram.na3_x1_49_ins.i0
* NET 887 = core.iram.na3_x1_16_sig
* NET 888 = core.iram.na3_x1_15_sig
* NET 892 = core.iram.a3_x2_5_sig
* NET 896 = core.iram.na3_x1_18_sig
* NET 898 = core.iram.a2_x2_5_sig
* NET 900 = core.iram.na3_x1_19_sig
* NET 903 = core.iram.na3_x1_19_ins.i0
* NET 904 = core.iram.ab_data_idx_1[1]
* NET 907 = core.iram.na3_x1_51_sig
* NET 908 = core.iram.na3_x1_49_sig
* NET 913 = core.iram.ab_data_idx_0[1]
* NET 914 = core.iram.na3_x1_50_sig
* NET 917 = core.iram.a2_x2_10_sig
* NET 921 = core.iram.na3_x1_48_sig
* NET 926 = core.iram.ab_data_idx_4[1]
* NET 929 = core.iram.no2_x1_15_sig
* NET 930 = core.iram.noa2a2a2a24_x1_3_sig
* NET 932 = core.iram.no2_x1_17_ins.i0
* NET 933 = core.iram.no2_x1_17_sig
* NET 934 = core.iram.na2_x1_28_sig
* NET 937 = core.iram.na2_x1_29_sig
* NET 938 = core.iram.ao22_x2_27_sig
* NET 941 = core.iram.ab_data_idx_6_1_ins.sff_s
* NET 943 = core.iram.ao22_x2_26_sig
* NET 944 = core.iram.ab_data_idx_6_1_ins.y
* NET 945 = core.iram.ab_data_idx_6_1_ins.sff_m
* NET 949 = core.iram.ab_data_idx_6_1_ins.u
* NET 950 = core.iram.ab_data_idx_6_1_ins.ckr
* NET 951 = core.iram.ab_data_idx_6_1_ins.nckr
* NET 952 = p_zero.137nymous_
* NET 988 = core.iram.aux157_ins.i0
* NET 993 = p_b0.639nymous_
* NET 994 = p_b0.132nymous_
* NET 995 = p_zero.69onymous_
* NET 996 = p_zero.74onymous_
* NET 1000 = core.iram.o2_x2_sig
* NET 1001 = core.iram.inv_x2_14_sig
* NET 1004 = core.iram.na4_x1_sig
* NET 1007 = core.iram.no2_x1_sig
* NET 1008 = core.iram.on12_x1_sig
* NET 1011 = core.iram.ab_data_idx_13_1_ins.y
* NET 1012 = core.iram.ab_data_idx_13_1_ins.sff_s
* NET 1013 = core.iram.oa2a2a23_x2_sig
* NET 1014 = core.iram.ab_data_idx_13_1_ins.ckr
* NET 1015 = core.iram.ab_data_idx_13_1_ins.u
* NET 1016 = core.iram.ab_data_idx_13_1_ins.sff_m
* NET 1020 = core.iram.ab_data_idx_13_1_ins.ck
* NET 1021 = core.iram.ab_data_idx_13_1_ins.nckr
* NET 1026 = core.iram.not_aux71_ins.i0
* NET 1027 = core.iram.no2_x1_12_ins.i0
* NET 1030 = core.iram.ab_data_idx_12[1]
* NET 1032 = core.iram.ab_data_idx_13[1]
* NET 1033 = core.iram.no2_x1_13_sig
* NET 1035 = core.iram.no2_x1_12_sig
* NET 1037 = core.iram.noa2a2a23_x1_sig
* NET 1040 = core.iram.not_aux71
* NET 1042 = core.iram.no2_x1_46_ins.i0
* NET 1044 = core.iram.ab_data_idx_15[1]
* NET 1045 = core.iram.no2_x1_46_sig
* NET 1049 = core.iram.no2_x1_45_sig
* NET 1051 = core.iram.ab_data_idx_11[1]
* NET 1053 = core.iram.noa2a2a23_x1_4_sig
* NET 1055 = core.iram.na2_x1_52_sig
* NET 1056 = core.iram.na3_x1_21_sig
* NET 1057 = core.iram.na4_x1_4_sig
* NET 1058 = core.iram.na4_x1_5_sig
* NET 1061 = core.iram.ab_data_idx_10[1]
* NET 1062 = core.iram.na3_x1_17_sig
* NET 1063 = core.iram.ab_data_idx_5[1]
* NET 1064 = core.iram.na3_x1_45_sig
* NET 1065 = core.iram.na3_x1_45_ins.i0
* NET 1066 = core.iram.na3_x1_20_sig
* NET 1067 = core.iram.a2_x2_9_sig
* NET 1068 = core.iram.a3_x2_10_sig
* NET 1069 = core.iram.a4_x2_2_sig
* NET 1070 = core.iram.na3_x1_22_sig
* NET 1072 = core.iram.na3_x1_20_ins.i0
* NET 1074 = core.iram.ab_data_idx_2_1_ins.sff_s
* NET 1075 = core.iram.ab_data_idx_2_1_ins.y
* NET 1077 = core.iram.ab_data_idx_2_1_ins.u
* NET 1078 = core.iram.ab_data_idx_2_1_ins.sff_m
* NET 1080 = core.iram.ab_data_idx_2_1_ins.ckr
* NET 1082 = core.iram.ao22_x2_10_sig
* NET 1083 = core.iram.ab_data_idx_2_1_ins.nckr
* NET 1084 = core.iram.na2_x1_12_sig
* NET 1088 = core.iram.no2_x1_16_sig
* NET 1090 = core.iram.ab_data_idx_3[1]
* NET 1091 = core.iram.ab_data_idx_2[1]
* NET 1092 = core.iram.ab_data_idx_6[1]
* NET 1095 = core.iram.ab_data_idx_7[1]
* NET 1096 = core.iram.noa2a2a2a24_x1_8_sig
* NET 1098 = core.iram.no2_x1_51_sig
* NET 1103 = core.iram.no2_x1_50_sig
* NET 1104 = p_b0.80onymous_
* NET 1105 = p_b0.57onymous_
* NET 1106 = p_zero.n16b
* NET 1111 = core.iram.not_aux138
* NET 1116 = core.iram.no4_x1_sig
* NET 1117 = core.iram.not_aux140_ins.i0
* NET 1123 = core.iram.o4_x2_sig
* NET 1126 = core.iram.not_b_2_ins.i
* NET 1128 = core.iram.ab_data_idx_14_1_ins.sff_s
* NET 1129 = core.iram.ab_data_idx_14_1_ins.y
* NET 1130 = core.iram.ab_data_idx_14_1_ins.sff_m
* NET 1133 = core.iram.na3_x1_4_sig
* NET 1134 = core.iram.ab_data_idx_14_1_ins.ck
* NET 1135 = core.iram.ab_data_idx_14_1_ins.u
* NET 1136 = core.iram.ab_data_idx_14_1_ins.ckr
* NET 1137 = core.iram.ab_data_idx_14_1_ins.nckr
* NET 1138 = core.iram.na2_x1_51_sig
* NET 1143 = core.iram.inv_x2_17_sig
* NET 1147 = core.iram.no2_x1_14_sig
* NET 1148 = core.iram.nao22_x1_6_ins.i0
* NET 1150 = core.iram.nao22_x1_6_sig
* NET 1152 = core.iram.ab_data_idx_8[2]
* NET 1156 = core.iram.a3_x2_13_sig
* NET 1159 = core.iram.a3_x2_11_ins.i0
* NET 1160 = core.iram.ab_data_idx_8[1]
* NET 1166 = core.iram.no2_x1_19_sig
* NET 1167 = core.iram.a3_x2_11_sig
* NET 1169 = core.iram.noa22_x1_8_sig
* NET 1170 = core.iram.ao22_x2_39_ins.i0
* NET 1175 = core.iram.na3_x1_54_sig
* NET 1176 = core.iram.na3_x1_53_sig
* NET 1179 = core.iram.a3_x2_6_sig
* NET 1180 = core.iram.o3_x2_6_sig
* NET 1184 = core.iram.noa22_x1_9_sig
* NET 1188 = core.iram.a4_x2_3_sig
* NET 1189 = core.iram.a3_x2_12_sig
* NET 1192 = core.iram.a2_x2_12_sig
* NET 1193 = core.iram.a2_x2_11_sig
* NET 1196 = core.iram.na3_x1_52_sig
* NET 1198 = core.iram.na3_x1_52_ins.i0
* NET 1200 = core.iram.na2_x1_25_sig
* NET 1204 = core.iram.no2_x1_21_ins.i0
* NET 1206 = core.iram.ab_data_idx_4[2]
* NET 1207 = core.iram.no2_x1_21_sig
* NET 1214 = core.iram.noa2a2a2a24_x1_4_sig
* NET 1216 = core.iram.no2_x1_22_sig
* NET 1219 = core.iram.no2_x1_20_sig
* NET 1221 = core.iram.no2_x1_49_sig
* NET 1225 = core.iram.no2_x1_57_sig
* NET 1226 = core.iram.ab_data_idx_6[2]
* NET 1231 = core.iram.no2_x1_58_sig
* NET 1232 = core.iram.ab_data_idx_7[2]
* NET 1235 = core.iram.noa2a2a2a24_x1_9_sig
* NET 1236 = core.iram.no2_x1_59_ins.i0
* NET 1238 = core.iram.no2_x1_59_sig
* NET 1239 = p_b0.1280ymous_
* NET 1240 = p_b0.cpb
* NET 1241 = p_b0.324nymous_
* NET 1243 = p_zero.p6c
* NET 1244 = p_zero.301nymous_
* NET 1245 = p_zero.305nymous_
* NET 1246 = p_zero.274nymous_
* NET 1278 = p_b0.259nymous_
* NET 1279 = p_zero.227nymous_
* NET 1280 = zero
* NET 1281 = p_zero.197nymous_
* NET 1282 = p_zero.224nymous_
* NET 1283 = p_zero.193nymous_
* NET 1284 = core.iram.not_aux20_ins.i1
* NET 1287 = core.iram.not_aux20
* NET 1288 = core.iram.o3_x2_2_sig
* NET 1294 = core.iram.not_aux21
* NET 1297 = core.iram.no3_x1_4_sig
* NET 1298 = core.iram.ab_data_idx_14[1]
* NET 1299 = core.iram.nao22_x1_5_sig
* NET 1302 = core.iram.not_aux30
* NET 1306 = core.iram.ab_data_idx_15_2_ins.sff_s
* NET 1307 = core.iram.ab_data_idx_15_2_ins.y
* NET 1308 = core.iram.ab_data_idx_15_2_ins.sff_m
* NET 1311 = core.iram.ao22_x2_50_sig
* NET 1312 = core.iram.ab_data_idx_15_2_ins.u
* NET 1313 = core.iram.ab_data_idx_15_2_ins.ckr
* NET 1315 = core.iram.not_aux80_ins.i0
* NET 1316 = core.iram.ab_data_idx_15_2_ins.nckr
* NET 1318 = core.iram.not_aux80_ins.i1
* NET 1323 = core.iram.no2_x1_24_ins.i0
* NET 1326 = core.iram.ab_data_idx_12[2]
* NET 1328 = core.iram.ab_data_idx_15[2]
* NET 1329 = core.iram.no2_x1_25_sig
* NET 1330 = core.iram.no2_x1_24_sig
* NET 1331 = core.iram.noa2a2a2a24_x1_5_sig
* NET 1337 = core.iram.no2_x1_27_sig
* NET 1338 = core.iram.no2_x1_47_sig
* NET 1339 = core.iram.no2_x1_52_sig
* NET 1343 = core.iram.no2_x1_54_sig
* NET 1345 = core.iram.noa2a2a23_x1_5_sig
* NET 1347 = core.iram.ab_data_idx_11[2]
* NET 1348 = core.iram.ab_data_idx_10[2]
* NET 1349 = core.iram.na3_x1_26_ins.i0
* NET 1350 = core.iram.na3_x1_26_sig
* NET 1351 = core.iram.na3_x1_28_sig
* NET 1352 = core.iram.na4_x1_6_sig
* NET 1353 = core.iram.na4_x1_7_sig
* NET 1357 = core.iram.ab_data_idx_5[2]
* NET 1358 = core.iram.ab_data_idx_5_2_ins.y
* NET 1360 = core.iram.ab_data_idx_5_2_ins.sff_m
* NET 1361 = core.iram.ab_data_idx_5_2_ins.sff_s
* NET 1362 = core.iram.ab_data_idx_5_2_ins.ck
* NET 1363 = core.iram.ao22_x2_23_sig
* NET 1364 = core.iram.ab_data_idx_5_2_ins.u
* NET 1366 = core.iram.ab_data_idx_5_2_ins.ckr
* NET 1367 = core.iram.ab_data_idx_5_2_ins.nckr
* NET 1368 = core.iram.na3_x1_29_sig
* NET 1369 = core.iram.no2_x1_23_sig
* NET 1371 = core.iram.ab_data_idx_3[2]
* NET 1372 = core.iram.na3_x1_27_sig
* NET 1373 = core.iram.no2_x1_48_ins.i0
* NET 1374 = core.iram.no2_x1_48_sig
* NET 1377 = core.iram.no2_x1_18_sig
* NET 1379 = core.iram.na2_x1_13_sig
* NET 1382 = core.iram.ab_data_idx_2[2]
* NET 1384 = core.iram.ab_data_idx_2_2_ins.sff_s
* NET 1385 = core.iram.ao22_x2_11_sig
* NET 1386 = core.iram.ab_data_idx_2_2_ins.y
* NET 1389 = core.iram.ab_data_idx_2_2_ins.sff_m
* NET 1392 = core.iram.ab_data_idx_2_2_ins.u
* NET 1393 = core.iram.ab_data_idx_2_2_ins.ckr
* NET 1394 = core.iram.ab_data_idx_2_2_ins.nckr
* NET 1396 = core.iram.no2_x1_56_sig
* NET 1398 = p_b0.1066ymous_
* NET 1400 = p_b0.n14c
* NET 1402 = b[0]
* NET 1403 = p_zero.318nymous_
* NET 1405 = core.iram.not_aux7_ins.i1
* NET 1407 = core.iram.not_alu_out[0]
* NET 1411 = core.iram.inv_x2_2_sig
* NET 1412 = core.iram.not_aux95
* NET 1413 = core.iram.not_aux8_ins.i0
* NET 1415 = core.iram.not_aux91_ins.i0
* NET 1421 = core.iram.aux154
* NET 1426 = core.iram.not_aux80
* NET 1428 = core.iram.aux81_ins.nq
* NET 1434 = core.iram.ab_data_idx_14_2_ins.ck
* NET 1435 = core.iram.ab_data_idx_14_2_ins.u
* NET 1436 = core.iram.ab_data_idx_14_2_ins.ckr
* NET 1437 = core.iram.ab_data_idx_14_2_ins.nckr
* NET 1438 = core.iram.na2_x1_48_sig
* NET 1440 = core.iram.ao22_x2_47_sig
* NET 1441 = core.iram.ab_data_idx_14[2]
* NET 1442 = core.iram.no2_x1_26_ins.i0
* NET 1445 = core.iram.no2_x1_26_sig
* NET 1449 = core.iram.no2_x1_44_sig
* NET 1451 = core.iram.no2_x1_55_sig
* NET 1452 = core.iram.no2_x1_53_ins.i0
* NET 1454 = core.iram.no2_x1_53_sig
* NET 1460 = core.iram.aux61_ins.i0
* NET 1465 = core.iram.aux14_ins.i0
* NET 1472 = core.iram.not_aux55
* NET 1474 = core.iram.na2_x1_27_sig
* NET 1478 = core.iram.ao22_x2_25_sig
* NET 1483 = core.iram.ab_data_idx_6_0_ins.u
* NET 1485 = core.iram.ab_data_idx_6_0_ins.ckr
* NET 1486 = core.iram.ab_data_idx_6_0_ins.nckr
* NET 1492 = core.iram.aux17
* NET 1499 = core.iram.na3_x1_3_ins.i1
* NET 1507 = core.iram.ab_data_idx_14_2_ins.sff_s
* NET 1509 = core.iram.ab_data_idx_14_2_ins.y
* NET 1510 = core.iram.ab_data_idx_14_2_ins.sff_m
* NET 1516 = core.iram.not_aux8
* NET 1522 = core.iram.aux159
* NET 1527 = core.iram.not_aux9
* NET 1532 = core.iram.aux160
* NET 1541 = core.iram.ab_data_idx_6_0_ins.sff_s
* NET 1542 = core.iram.ab_data_idx_6_0_ins.sff_m
* NET 1543 = core.iram.ab_data_idx_6_0_ins.y
* NET 1548 = p_a3.132nymous_
* NET 1549 = p_ovr.n15d
* NET 1550 = p_ovr.n18f
* NET 1551 = core.iram.not_aux101_ins.i0
* NET 1552 = core.iram.not_aux15
* NET 1560 = core.iram.r0_to_ins.q
* NET 1563 = core.iram.no2_x1_68_sig
* NET 1564 = core.iram.not_b[0]
* NET 1565 = core.iram.not_aux7
* NET 1569 = core.iram.not_aux43
* NET 1575 = core.iram.ab_data_idx_15_0_ins.y
* NET 1576 = core.iram.ab_data_idx_15_0_ins.sff_s
* NET 1577 = core.iram.ab_data_idx_15_0_ins.u
* NET 1579 = core.iram.ab_data_idx_15_0_ins.sff_m
* NET 1581 = core.iram.ab_data_idx_15_0_ins.ck
* NET 1582 = core.iram.ao22_x2_49_sig
* NET 1583 = core.iram.ab_data_idx_15_0_ins.ckr
* NET 1584 = core.iram.ab_data_idx_15_0_ins.nckr
* NET 1585 = core.iram.aux103
* NET 1588 = core.iram.na2_x1_50_sig
* NET 1589 = core.iram.not_aux69
* NET 1591 = core.iram.not_b[3]
* NET 1592 = core.iram.not_aux46_ins.i0
* NET 1595 = core.iram.aux87_ins.i0
* NET 1598 = core.iram.not_aux46
* NET 1600 = core.iram.na2_x1_39_sig
* NET 1604 = core.iram.ab_data_idx_10_0_ins.y
* NET 1606 = core.iram.ab_data_idx_10_0_ins.sff_m
* NET 1607 = core.iram.ab_data_idx_10_0_ins.sff_s
* NET 1608 = core.iram.ao22_x2_37_sig
* NET 1610 = core.iram.ab_data_idx_10_0_ins.u
* NET 1612 = core.iram.ab_data_idx_10_0_ins.ckr
* NET 1613 = core.iram.ab_data_idx_10_0_ins.nckr
* NET 1615 = core.iram.ab_data_idx_0_0_ins.y
* NET 1617 = core.iram.ab_data_idx_0_0_ins.sff_s
* NET 1618 = core.iram.ab_data_idx_0_0_ins.u
* NET 1620 = core.iram.ab_data_idx_0_0_ins.sff_m
* NET 1621 = core.iram.ab_data_idx_0_0_ins.ckr
* NET 1622 = core.iram.ab_data_idx_0_0_ins.ck
* NET 1623 = core.iram.ab_data_idx_0_0_ins.nckr
* NET 1624 = core.iram.ao22_x2_sig
* NET 1627 = core.iram.na2_x1_3_sig
* NET 1628 = core.iram.ab_data_idx_3_0_ins.y
* NET 1630 = core.iram.ab_data_idx_3_0_ins.sff_s
* NET 1631 = core.iram.ab_data_idx_3_0_ins.ckr
* NET 1632 = core.iram.ab_data_idx_3_0_ins.u
* NET 1635 = core.iram.ab_data_idx_3_0_ins.sff_m
* NET 1637 = core.iram.ab_data_idx_3_0_ins.nckr
* NET 1638 = core.iram.ao22_x2_13_sig
* NET 1641 = core.iram.na2_x1_15_sig
* NET 1642 = core.iram.na2_x1_11_sig
* NET 1646 = core.iram.not_aux115
* NET 1650 = core.iram.ab_data_idx_2_0_ins.sff_s
* NET 1651 = core.iram.ao22_x2_9_sig
* NET 1652 = core.iram.ab_data_idx_2_0_ins.y
* NET 1654 = core.iram.ab_data_idx_2_0_ins.sff_m
* NET 1656 = core.iram.ab_data_idx_2_0_ins.ck
* NET 1657 = core.iram.ab_data_idx_2_0_ins.u
* NET 1658 = core.iram.ab_data_idx_2_0_ins.nckr
* NET 1659 = core.iram.ab_data_idx_2_0_ins.ckr
* NET 1660 = p_a3.93onymous_
* NET 1661 = p_a3.p2
* NET 1662 = p_ovr.406nymous_
* NET 1663 = p_ovr.13onymous_
* NET 1689 = p_a3.cpb
* NET 1690 = p_a3.414nymous_
* NET 1691 = p_a3.n8b
* NET 1693 = p_ovr.299nymous_
* NET 1694 = p_ovr.p7a
* NET 1695 = p_ovr.293nymous_
* NET 1696 = r0_from_pads
* NET 1697 = core.iram.na2_x1_2_sig
* NET 1700 = core.iram.a3_x2_ins.i2
* NET 1702 = core.iram.a3_x2_sig
* NET 1704 = core.iram.not_aux29
* NET 1706 = core.iram.na2_x1_sig
* NET 1708 = core.iram.inv_x2_4_sig
* NET 1710 = core.iram.not_aux78
* NET 1713 = core.iram.not_aux79_ins.i0
* NET 1716 = core.iram.ab_data_idx_9_0_ins.sff_s
* NET 1718 = core.iram.noa2a22_x1_sig
* NET 1719 = core.iram.ab_data_idx_9_0_ins.y
* NET 1722 = core.iram.ab_data_idx_9_0_ins.u
* NET 1723 = core.iram.ab_data_idx_9_0_ins.sff_m
* NET 1727 = core.iram.ab_data_idx_9_0_ins.ckr
* NET 1728 = core.iram.ab_data_idx_9_0_ins.nckr
* NET 1730 = core.iram.not_aux89
* NET 1736 = core.iram.ab_data_idx_11_0_ins.y
* NET 1737 = core.iram.ab_data_idx_11_0_ins.sff_s
* NET 1738 = core.iram.noa2a22_x1_2_sig
* NET 1739 = core.iram.ab_data_idx_11_0_ins.u
* NET 1741 = core.iram.ab_data_idx_11_0_ins.sff_m
* NET 1743 = core.iram.ab_data_idx_11_0_ins.ckr
* NET 1744 = core.iram.ab_data_idx_11_0_ins.ck
* NET 1745 = core.iram.ab_data_idx_11_0_ins.nckr
* NET 1747 = core.iram.inv_x2_8_sig
* NET 1750 = core.iram.not_aux85
* NET 1751 = core.iram.na2_x1_47_sig
* NET 1754 = core.iram.aux155
* NET 1755 = core.iram.aux102_ins.i0
* NET 1764 = core.iram.na3_x1_40_sig
* NET 1765 = core.iram.na3_x1_39_sig
* NET 1770 = core.iram.no2_x1_38_ins.i0
* NET 1782 = core.iram.not_aux60_ins.i1
* NET 1785 = core.iram.not_aux44
* NET 1789 = core.iram.na3_x1_13_sig
* NET 1790 = core.iram.na3_x1_11_sig
* NET 1794 = core.iram.na3_x1_12_ins.i0
* NET 1797 = core.iram.na3_x1_12_sig
* NET 1798 = core.iram.a2_x2_8_sig
* NET 1804 = core.iram.not_aux60
* NET 1809 = core.iram.na3_x1_14_sig
* NET 1810 = core.iram.ab_data_idx_3[0]
* NET 1812 = core.iram.ab_data_idx_2[0]
* NET 1813 = core.iram.no2_x1_41_sig
* NET 1815 = core.iram.noa2a2a2a24_x1_7_sig
* NET 1819 = core.iram.no2_x1_43_sig
* NET 1821 = core.iram.no2_x1_40_sig
* NET 1825 = core.iram.no2_x1_42_sig
* NET 1826 = p_a3.259nymous_
* NET 1827 = p_a3.1280ymous_
* NET 1828 = ovr
* NET 1829 = p_ovr.p3
* NET 1830 = p_ovr.n3
* NET 1831 = p_ovr.224nymous_
* NET 1834 = core.iram.na3_x1_ins.i1
* NET 1838 = core.iram.not_aux142
* NET 1842 = core.iram.na3_x1_ins.i0
* NET 1843 = core.iram.na3_x1_sig
* NET 1844 = core.iram.aux4_ins.i1
* NET 1847 = core.iram.aux4
* NET 1849 = core.iram.not_aux116_ins.i1
* NET 1852 = core.iram.ab_data_idx_12_0_ins.sff_s
* NET 1854 = core.iram.ab_data_idx_12_0_ins.y
* NET 1856 = core.iram.ab_data_idx_12_0_ins.u
* NET 1857 = core.iram.ab_data_idx_12_0_ins.sff_m
* NET 1860 = core.iram.ab_data_idx_12_0_ins.ckr
* NET 1861 = core.iram.ab_data_idx_12_0_ins.nckr
* NET 1862 = core.iram.not_aux70
* NET 1863 = core.iram.na2_x1_43_sig
* NET 1865 = core.iram.ao22_x2_41_sig
* NET 1868 = core.iram.ab_data_idx_14_0_ins.y
* NET 1869 = core.iram.ab_data_idx_14_0_ins.sff_s
* NET 1870 = core.iram.ao22_x2_46_sig
* NET 1872 = core.iram.ab_data_idx_14_0_ins.u
* NET 1874 = core.iram.ab_data_idx_14_0_ins.sff_m
* NET 1875 = core.iram.ab_data_idx_14_0_ins.ck
* NET 1876 = core.iram.ab_data_idx_14_0_ins.nckr
* NET 1877 = core.iram.ab_data_idx_14_0_ins.ckr
* NET 1878 = core.iram.ab_data_idx_9[0]
* NET 1879 = core.iram.na3_x1_9_ins.i0
* NET 1881 = core.iram.no2_x1_63_ins.i0
* NET 1882 = core.iram.not_aux109
* NET 1884 = core.iram.no2_x1_39_sig
* NET 1885 = core.iram.ab_data_idx_11[0]
* NET 1886 = core.iram.ab_data_idx_10[0]
* NET 1887 = core.iram.no2_x1_38_sig
* NET 1891 = core.iram.no2_x1_37_sig
* NET 1893 = core.iram.na3_x1_58_ins.i2
* NET 1894 = core.iram.not_aux116
* NET 1895 = core.iram.not_aux45
* NET 1896 = core.iram.not_aux10
* NET 1897 = core.iram.na2_x1_23_sig
* NET 1902 = core.iram.ab_data_idx_5_0_ins.sff_s
* NET 1903 = core.iram.ab_data_idx_5_0_ins.y
* NET 1905 = core.iram.ab_data_idx_5_0_ins.sff_m
* NET 1906 = core.iram.ao22_x2_21_sig
* NET 1908 = core.iram.ab_data_idx_5_0_ins.u
* NET 1909 = core.iram.ab_data_idx_5_0_ins.nckr
* NET 1910 = core.iram.ab_data_idx_5_0_ins.ckr
* NET 1911 = core.iram.na3_x1_12_ins.i2
* NET 1914 = core.iram.no2_x1_5_sig
* NET 1915 = core.iram.ab_data_idx_6[0]
* NET 1919 = core.iram.no2_x1_7_ins.i0
* NET 1920 = core.iram.no2_x1_7_sig
* NET 1923 = core.iram.no2_x1_4_sig
* NET 1925 = core.iram.na2_x1_31_sig
* NET 1928 = core.iram.ab_data_idx_7[0]
* NET 1930 = core.iram.ab_data_idx_7_0_ins.sff_s
* NET 1931 = core.iram.ao22_x2_29_sig
* NET 1932 = core.iram.ab_data_idx_7_0_ins.y
* NET 1935 = core.iram.ab_data_idx_7_0_ins.sff_m
* NET 1936 = core.iram.ab_data_idx_7_0_ins.ck
* NET 1937 = core.iram.ab_data_idx_7_0_ins.nckr
* NET 1938 = core.iram.ab_data_idx_7_0_ins.ckr
* NET 1939 = core.iram.ab_data_idx_7_0_ins.u
* NET 1940 = p_a3.196nymous_
* NET 1941 = a[3]
* NET 1942 = p_ovr.889nymous_
* NET 1943 = p_ovr.793nymous_
* NET 1970 = p_a3.n14a
* NET 1971 = p_a3.568nymous_
* NET 1972 = core.iram.not_i[2]
* NET 1975 = core.iram.not_aux140
* NET 1976 = core.iram.not_aux101
* NET 1977 = core.iram.no3_x1_5_sig
* NET 1984 = core.iram.o3_x2_4_sig
* NET 1985 = core.iram.nao22_x1_8_sig
* NET 1988 = core.iram.ab_data_idx_13_0_ins.sff_s
* NET 1990 = core.iram.ab_data_idx_13_0_ins.y
* NET 1993 = core.iram.ab_data_idx_13_0_ins.sff_m
* NET 1996 = core.iram.ab_data_idx_13_0_ins.ckr
* NET 1997 = core.iram.ab_data_idx_13_0_ins.nckr
* NET 1998 = core.iram.ab_data_idx_13_0_ins.u
* NET 1999 = core.iram.aux153
* NET 2001 = core.iram.noa2ao222_x1_ins.i3
* NET 2002 = core.iram.not_aux124
* NET 2003 = core.iram.inv_x2_13_sig
* NET 2004 = core.iram.not_aux79
* NET 2005 = core.iram.noa2ao222_x1_sig
* NET 2008 = core.iram.inv_x2_12_sig
* NET 2012 = core.iram.na2_x1_35_sig
* NET 2020 = core.iram.aux156
* NET 2023 = core.iram.ab_data_idx_14[0]
* NET 2026 = core.iram.no2_x1_8_sig
* NET 2027 = core.iram.ab_data_idx_12[0]
* NET 2031 = core.iram.no2_x1_9_sig
* NET 2032 = core.iram.no2_x1_10_ins.i0
* NET 2033 = core.iram.no2_x1_10_sig
* NET 2034 = core.iram.na3_x1_40_ins.i2
* NET 2035 = core.iram.na3_x1_9_sig
* NET 2041 = core.iram.o3_x2_5_sig
* NET 2042 = core.iram.noa2a2a2a24_x1_sig
* NET 2043 = core.iram.a3_x2_4_sig
* NET 2044 = core.iram.noa2a2a2a24_x1_2_sig
* NET 2050 = core.iram.noa2a2a23_x1_3_sig
* NET 2055 = core.iram.ab_data_idx_13[0]
* NET 2064 = core.iram.na3_x1_10_sig
* NET 2065 = core.iram.ab_data_idx_5[0]
* NET 2066 = core.iram.na3_x1_38_sig
* NET 2070 = core.iram.ab_data_idx_0[0]
* NET 2075 = core.iram.na3_x1_42_sig
* NET 2076 = core.iram.na3_x1_43_sig
* NET 2081 = core.iram.na3_x1_41_ins.i0
* NET 2084 = core.iram.na3_x1_41_sig
* NET 2087 = core.iram.a2_x2_7_sig
* NET 2088 = core.iram.a3_x2_8_sig
* NET 2091 = core.iram.no2_x1_6_ins.i0
* NET 2092 = core.iram.a4_x2_sig
* NET 2094 = core.iram.no2_x1_6_sig
* NET 2096 = core.iram.na2_x1_19_sig
* NET 2099 = core.iram.ab_data_idx_4[0]
* NET 2101 = core.iram.ab_data_idx_4_0_ins.y
* NET 2103 = core.iram.ab_data_idx_4_0_ins.sff_m
* NET 2104 = core.iram.ab_data_idx_4_0_ins.sff_s
* NET 2105 = core.iram.ab_data_idx_4_0_ins.ck
* NET 2106 = core.iram.ao22_x2_17_sig
* NET 2107 = core.iram.ab_data_idx_4_0_ins.u
* NET 2108 = core.iram.ab_data_idx_4_0_ins.ckr
* NET 2112 = core.iram.ab_data_idx_4_0_ins.nckr
* NET 2118 = core.iram.aux158
* NET 2121 = p_vddick0.267nymous_
* NET 2122 = core.iram.not_aux36_ins.i1
* NET 2126 = core.iram.ab_data_idx_15_3_ins.sff_m
* NET 2128 = core.iram.ab_data_idx_15_3_ins.sff_s
* NET 2129 = core.iram.ab_data_idx_15_3_ins.y
* NET 2130 = core.iram.na3_x1_7_sig
* NET 2132 = core.iram.ab_data_idx_15_3_ins.u
* NET 2134 = core.iram.ab_data_idx_15_3_ins.ckr
* NET 2135 = core.iram.ab_data_idx_15_3_ins.nckr
* NET 2136 = core.iram.not_alu_out[1]
* NET 2138 = core.iram.not_aux0
* NET 2140 = core.iram.inv_x2_15_sig
* NET 2143 = core.iram.na3_x1_3_sig
* NET 2146 = core.iram.o3_x2_3_ins.i1
* NET 2147 = core.iram.ao22_x2_45_sig
* NET 2149 = core.iram.ab_data_idx_8_0_ins.y
* NET 2151 = core.iram.ab_data_idx_8_0_ins.sff_s
* NET 2153 = core.iram.ao22_x2_33_sig
* NET 2154 = core.iram.ab_data_idx_8_0_ins.ckr
* NET 2155 = core.iram.ab_data_idx_8_0_ins.u
* NET 2157 = core.iram.ab_data_idx_8_0_ins.sff_m
* NET 2158 = core.iram.ab_data_idx_8_0_ins.ck
* NET 2159 = core.iram.ab_data_idx_8_0_ins.nckr
* NET 2160 = core.iram.inv_x2_16_sig
* NET 2161 = core.iram.ab_data_idx_8[0]
* NET 2165 = core.iram.no2_x1_11_sig
* NET 2167 = core.iram.a3_x2_9_sig
* NET 2168 = core.iram.ab_data_idx_15[0]
* NET 2170 = core.iram.noa22_x1_7_sig
* NET 2171 = core.iram.not_aux86
* NET 2173 = core.iram.no2_x1_36_sig
* NET 2175 = core.iram.not_aux111
* NET 2176 = core.iram.no2_x1_62_ins.i0
* NET 2178 = core.iram.na3_x1_8_ins.i0
* NET 2179 = core.iram.na3_x1_8_sig
* NET 2180 = core.iram.ab_data_idx_1_0_ins.y
* NET 2183 = core.iram.ab_data_idx_1_0_ins.sff_s
* NET 2184 = core.iram.ab_data_idx_1_0_ins.ckr
* NET 2185 = core.iram.ab_data_idx_1_0_ins.u
* NET 2187 = core.iram.ab_data_idx_1_0_ins.sff_m
* NET 2189 = core.iram.ao22_x2_5_sig
* NET 2190 = core.iram.ab_data_idx_1_0_ins.nckr
* NET 2191 = core.iram.na2_x1_7_sig
* NET 2195 = core.iram.ab_data_idx_1[0]
* NET 2196 = core.iram.na3_x1_44_sig
* NET 2197 = core.iram.aux12
* NET 2199 = core.iram.aux66
* NET 2202 = core.iram.na4_x1_3_sig
* NET 2203 = core.iram.na4_x1_2_sig
* NET 2208 = core.iram.ab_data_idx_0_3_ins.sff_s
* NET 2209 = core.iram.ab_data_idx_0_3_ins.y
* NET 2210 = core.iram.ab_data_idx_0_3_ins.ckr
* NET 2211 = core.iram.ab_data_idx_0_3_ins.u
* NET 2213 = core.iram.ab_data_idx_0_3_ins.sff_m
* NET 2214 = core.iram.ab_data_idx_0_3_ins.ck
* NET 2215 = core.iram.ao22_x2_4_sig
* NET 2216 = core.iram.ab_data_idx_0_3_ins.nckr
* NET 2217 = core.iram.aux14
* NET 2220 = core.iram.not_aux56
* NET 2222 = core.iram.not_aux61
* NET 2223 = core.iram.no2_x1_31_ins.i0
* NET 2226 = core.iram.no2_x1_67_ins.i0
* NET 2227 = core.iram.aux62
* NET 2229 = core.iram.not_aux114
* NET 2232 = core.iram.ab_data_idx_3_3_ins.sff_s
* NET 2233 = core.iram.ao22_x2_16_sig
* NET 2234 = core.iram.ab_data_idx_3_3_ins.y
* NET 2237 = core.iram.ab_data_idx_3_3_ins.sff_m
* NET 2239 = core.iram.ab_data_idx_3_3_ins.u
* NET 2240 = core.iram.ab_data_idx_3_3_ins.nckr
* NET 2241 = core.iram.ab_data_idx_3_3_ins.ckr
* NET 2242 = p_a2.112nymous_
* NET 2243 = p_a2.640nymous_
* NET 2282 = p_a2.43onymous_
* NET 2283 = p_a2.466nymous_
* NET 2284 = core.iram.not_alu_out[2]
* NET 2285 = core.iram.o3_x2_sig
* NET 2290 = core.iram.not_aux38
* NET 2295 = core.iram.nao22_x1_9_sig
* NET 2297 = core.iram.not_aux82
* NET 2301 = core.iram.no3_x1_sig
* NET 2303 = core.iram.ab_data_idx_11_3_ins.y
* NET 2305 = core.iram.ab_data_idx_11_3_ins.sff_s
* NET 2308 = core.iram.ab_data_idx_11_3_ins.u
* NET 2309 = core.iram.ab_data_idx_11_3_ins.ckr
* NET 2311 = core.iram.ab_data_idx_11_3_ins.sff_m
* NET 2312 = core.iram.ab_data_idx_11_3_ins.ck
* NET 2313 = core.iram.ab_data_idx_11_3_ins.nckr
* NET 2315 = core.iram.not_aux91
* NET 2317 = core.iram.noa22_x1_4_sig
* NET 2320 = core.iram.inv_x2_11_sig
* NET 2322 = core.iram.no3_x1_2_sig
* NET 2323 = core.iram.aux120
* NET 2324 = core.iram.no2_x1_28_ins.i0
* NET 2325 = core.iram.not_aux90
* NET 2327 = core.iram.no2_x1_28_sig
* NET 2328 = core.iram.no2_x1_29_sig
* NET 2332 = core.iram.no2_x1_30_sig
* NET 2335 = core.iram.not_aux105
* NET 2337 = core.iram.not_aux107
* NET 2341 = core.iram.no2_x1_63_sig
* NET 2345 = core.iram.no2_x1_62_sig
* NET 2346 = core.iram.no2_x1_61_sig
* NET 2355 = core.iram.na3_x1_36_ins.i0
* NET 2356 = core.iram.ab_data_idx_11[3]
* NET 2357 = core.iram.aux90
* NET 2360 = core.iram.aux48
* NET 2366 = core.iram.na2_x1_10_sig
* NET 2370 = core.iram.ab_data_idx_5_3_ins.sff_s
* NET 2372 = core.iram.ao22_x2_24_sig
* NET 2373 = core.iram.ab_data_idx_5_3_ins.y
* NET 2374 = core.iram.ab_data_idx_5_3_ins.u
* NET 2377 = core.iram.ab_data_idx_5_3_ins.sff_m
* NET 2379 = core.iram.ab_data_idx_5_3_ins.ckr
* NET 2380 = core.iram.ab_data_idx_5_3_ins.nckr
* NET 2384 = core.iram.no2_x1_33_sig
* NET 2388 = core.iram.no2_x1_31_sig
* NET 2390 = core.iram.not_aux12
* NET 2392 = core.iram.no2_x1_32_sig
* NET 2394 = core.iram.no2_x1_34_sig
* NET 2395 = core.iram.no2_x1_34_ins.i0
* NET 2399 = core.iram.na2_x1_6_sig
* NET 2401 = core.iram.na2_x1_18_sig
* NET 2402 = core.iram.no2_x1_67_sig
* NET 2404 = core.iram.no2_x1_65_sig
* NET 2410 = core.iram.not_aux112
* NET 2411 = core.iram.no2_x1_64_sig
* NET 2414 = core.iram.not_aux113
* NET 2415 = core.iram.no2_x1_66_ins.i0
* NET 2416 = core.iram.no2_x1_66_sig
* NET 2417 = p_a2.n6a
* NET 2418 = p_a2.1280ymous_
* NET 2419 = p_a2.n8a
* NET 2420 = p_a2.324nymous_
* NET 2421 = p_vddick0.14onymous_
* NET 2422 = p_vddick0.5nonymous_
* NET 2423 = core.iram.not_b[2]
* NET 2424 = core.iram.not_aux41
* NET 2426 = core.iram.inv_x2_7_sig
* NET 2427 = core.iram.ab_data_idx_13_2_ins.ck
* NET 2429 = core.iram.aux73
* NET 2432 = core.iram.na2_x1_38_sig
* NET 2435 = core.iram.aux72
* NET 2439 = core.iram.na3_x1_32_sig
* NET 2440 = core.iram.na3_x1_31_sig
* NET 2443 = core.iram.noa2a2a2a24_x1_6_sig
* NET 2444 = core.iram.noa2a2a23_x1_2_sig
* NET 2445 = core.iram.na3_x1_33_sig
* NET 2447 = core.iram.aux47
* NET 2448 = core.iram.na3_x1_34_ins.i0
* NET 2449 = core.iram.na3_x1_34_sig
* NET 2450 = core.iram.na3_x1_30_sig
* NET 2451 = core.iram.ab_data_idx_1_3_ins.ck
* NET 2453 = core.iram.na2_x1_26_sig
* NET 2455 = core.iram.aux65
* NET 2457 = core.iram.not_aux147
* NET 2459 = core.iram.na2_x1_22_sig
* NET 2462 = core.iram.na2_x1_34_sig
* NET 2465 = core.iram.ab_data_idx_7_3_ins.ck
* NET 2466 = p_a2.nnt
* NET 2467 = a[2]
* NET 2468 = core.iram.no2_x1_2_ins.i0
* NET 2471 = core.iram.no3_x1_3_ins.i2
* NET 2472 = core.iram.o2_x2_4_sig
* NET 2476 = core.iram.o2_x2_3_sig
* NET 2479 = core.iram.no3_x1_3_sig
* NET 2483 = core.iram.noa22_x1_6_sig
* NET 2485 = core.iram.ab_data_idx_13_2_ins.ckr
* NET 2486 = core.iram.ab_data_idx_13_2_ins.nckr
* NET 2487 = core.iram.ab_data_idx_13_2_ins.sff_m
* NET 2488 = core.iram.ab_data_idx_13[2]
* NET 2490 = core.iram.ab_data_idx_13_2_ins.sff_s
* NET 2491 = core.iram.ab_data_idx_13_2_ins.y
* NET 2494 = core.iram.ab_data_idx_13_2_ins.u
* NET 2497 = core.iram.ab_data_idx_8[3]
* NET 2498 = core.iram.ab_data_idx_8_3_ins.ckr
* NET 2499 = core.iram.ab_data_idx_8_3_ins.nckr
* NET 2500 = core.iram.ab_data_idx_8_3_ins.sff_m
* NET 2502 = core.iram.ab_data_idx_8_3_ins.sff_s
* NET 2503 = core.iram.ab_data_idx_8_3_ins.y
* NET 2507 = core.iram.ab_data_idx_8_3_ins.u
* NET 2511 = core.iram.ao22_x2_36_sig
* NET 2513 = core.iram.not_aux72
* NET 2516 = core.iram.ab_data_idx_15[3]
* NET 2517 = core.iram.no2_x1_60_sig
* NET 2520 = core.iram.a3_x2_15_sig
* NET 2526 = core.iram.a3_x2_7_sig
* NET 2529 = core.iram.a2_x2_6_sig
* NET 2532 = core.iram.ab_data_idx_1_3_ins.ckr
* NET 2533 = core.iram.ab_data_idx_1_3_ins.nckr
* NET 2534 = core.iram.ab_data_idx_1_3_ins.sff_m
* NET 2535 = core.iram.ab_data_idx_1_3_ins.sff_s
* NET 2537 = core.iram.ab_data_idx_1_3_ins.y
* NET 2538 = core.iram.ao22_x2_8_sig
* NET 2541 = core.iram.ab_data_idx_1_3_ins.u
* NET 2542 = core.iram.not_aux47
* NET 2544 = core.iram.not_aux148
* NET 2546 = core.iram.ab_data_idx_4_3_ins.ckr
* NET 2548 = core.iram.ab_data_idx_4_3_ins.nckr
* NET 2549 = core.iram.ab_data_idx_4_3_ins.sff_m
* NET 2551 = core.iram.ab_data_idx_4_3_ins.y
* NET 2552 = core.iram.ab_data_idx_4_3_ins.sff_s
* NET 2554 = core.iram.ab_data_idx_4_3_ins.u
* NET 2556 = core.iram.ao22_x2_20_sig
* NET 2559 = core.iram.ab_data_idx_7_3_ins.ckr
* NET 2560 = core.iram.ab_data_idx_7_3_ins.nckr
* NET 2561 = core.iram.ab_data_idx_7[3]
* NET 2562 = core.iram.ab_data_idx_7_3_ins.sff_s
* NET 2565 = core.iram.ab_data_idx_7_3_ins.y
* NET 2566 = core.iram.ao22_x2_32_sig
* NET 2567 = core.iram.ab_data_idx_7_3_ins.sff_m
* NET 2572 = core.iram.ab_data_idx_7_3_ins.u
* NET 2573 = p_a2.nt
* NET 2574 = p_a2.n14b
* NET 2575 = p_a2.87onymous_
* NET 2577 = core.iram.no2_x1_2_sig
* NET 2581 = core.iram.oa2ao222_x2_sig
* NET 2582 = core.iram.noa22_x1_5_sig
* NET 2584 = core.iram.not_aux36
* NET 2585 = core.iram.no2_x1_3_ins.i0
* NET 2586 = core.iram.no2_x1_3_sig
* NET 2587 = core.iram.o2_x2_2_sig
* NET 2592 = core.iram.o3_x2_3_sig
* NET 2593 = core.iram.a2_x2_sig
* NET 2594 = core.iram.nao22_x1_sig
* NET 2596 = core.iram.na3_x1_2_sig
* NET 2600 = core.iram.not_ab_data_idx_13[2]
* NET 2601 = core.iram.nao22_x1_2_sig
* NET 2604 = core.iram.ab_data_idx_12_3_ins.sff_s
* NET 2605 = core.iram.ab_data_idx_12_3_ins.y
* NET 2607 = core.iram.ab_data_idx_12_3_ins.sff_m
* NET 2610 = core.iram.ab_data_idx_12_3_ins.ckr
* NET 2611 = core.iram.ab_data_idx_12_3_ins.nckr
* NET 2612 = core.iram.ab_data_idx_12_3_ins.u
* NET 2613 = core.iram.aux93
* NET 2614 = core.iram.ao22_x2_44_sig
* NET 2617 = core.iram.not_aux151
* NET 2619 = core.iram.na2_x1_46_sig
* NET 2620 = core.iram.not_aux81
* NET 2621 = core.iram.no2_x1_35_ins.i0
* NET 2622 = core.iram.no2_x1_35_sig
* NET 2625 = core.iram.ab_data_idx_14_3_ins.y
* NET 2626 = core.iram.ab_data_idx_14_3_ins.sff_s
* NET 2628 = core.iram.ab_data_idx_14_3_ins.sff_m
* NET 2629 = core.iram.ab_data_idx_14_3_ins.ck
* NET 2630 = core.iram.ab_data_idx_14_3_ins.nckr
* NET 2631 = core.iram.ab_data_idx_14_3_ins.u
* NET 2633 = core.iram.ab_data_idx_14_3_ins.ckr
* NET 2634 = core.iram.ao22_x2_48_sig
* NET 2635 = core.iram.aux102
* NET 2636 = core.iram.ab_data_idx_14[3]
* NET 2639 = core.iram.na2_x1_49_sig
* NET 2641 = core.iram.na2_x1_42_sig
* NET 2643 = core.iram.ab_data_idx_10[3]
* NET 2645 = core.iram.ab_data_idx_10_3_ins.y
* NET 2646 = core.iram.ab_data_idx_10_3_ins.sff_s
* NET 2647 = core.iram.ao22_x2_40_sig
* NET 2648 = core.iram.ab_data_idx_10_3_ins.ckr
* NET 2649 = core.iram.ab_data_idx_10_3_ins.u
* NET 2651 = core.iram.ab_data_idx_10_3_ins.sff_m
* NET 2654 = core.iram.ab_data_idx_10_3_ins.nckr
* NET 2655 = core.iram.not_aux152
* NET 2656 = core.iram.aux86
* NET 2659 = core.iram.noa2a2a23_x1_6_sig
* NET 2660 = core.iram.noa22_x1_10_sig
* NET 2664 = core.iram.ab_data_idx_5[3]
* NET 2665 = core.iram.na3_x1_59_sig
* NET 2668 = core.iram.na4_x1_8_sig
* NET 2670 = core.iram.na3_x1_36_sig
* NET 2671 = core.iram.na3_x1_37_sig
* NET 2672 = core.iram.na2_x1_53_sig
* NET 2676 = core.iram.na4_x1_9_sig
* NET 2677 = core.iram.ab_data_idx_3[3]
* NET 2680 = core.iram.na3_x1_35_sig
* NET 2684 = core.iram.ab_data_idx_4[3]
* NET 2687 = core.iram.na3_x1_64_ins.i0
* NET 2688 = core.iram.ab_data_idx_0[3]
* NET 2694 = core.iram.not_aux150
* NET 2695 = core.iram.not_aux42
* NET 2696 = core.iram.aux56
* NET 2699 = core.iram.not_aux120
* NET 2701 = core.iram.na2_x1_14_sig
* NET 2702 = core.iram.aux57
* NET 2705 = core.iram.ab_data_idx_2[3]
* NET 2706 = core.iram.ab_data_idx_2_3_ins.sff_s
* NET 2708 = core.iram.ao22_x2_12_sig
* NET 2709 = core.iram.ab_data_idx_2_3_ins.y
* NET 2710 = core.iram.ab_data_idx_2_3_ins.sff_m
* NET 2713 = core.iram.ab_data_idx_2_3_ins.ck
* NET 2714 = core.iram.ab_data_idx_2_3_ins.u
* NET 2715 = core.iram.ab_data_idx_2_3_ins.ckr
* NET 2716 = core.iram.ab_data_idx_2_3_ins.nckr
* NET 2717 = p_np.137nymous_
* NET 2751 = p_a1.639nymous_
* NET 2752 = p_a1.132nymous_
* NET 2753 = p_np.69onymous_
* NET 2754 = p_np.74onymous_
* NET 2756 = core.iram.ab_data_idx_13_3_ins.sff_s
* NET 2757 = core.iram.ab_data_idx_13_3_ins.y
* NET 2759 = core.iram.ab_data_idx_13_3_ins.sff_m
* NET 2761 = core.iram.nao22_x1_4_sig
* NET 2762 = core.iram.ab_data_idx_13_3_ins.nckr
* NET 2763 = core.iram.ab_data_idx_13_3_ins.u
* NET 2765 = core.iram.ab_data_idx_13_3_ins.ckr
* NET 2766 = core.iram.not_i_1_ins.i
* NET 2768 = core.iram.ab_data_idx_9_3_ins.sff_m
* NET 2771 = core.iram.ab_data_idx_9_3_ins.sff_s
* NET 2772 = core.iram.ab_data_idx_9_3_ins.y
* NET 2773 = core.iram.ab_data_idx_9_3_ins.ck
* NET 2774 = core.iram.noa22_x1_3_sig
* NET 2775 = core.iram.ab_data_idx_9_3_ins.u
* NET 2776 = core.iram.ab_data_idx_9_3_ins.ckr
* NET 2777 = core.iram.ab_data_idx_9_3_ins.nckr
* NET 2778 = core.iram.not_alu_out[3]
* NET 2781 = core.iram.aux42
* NET 2782 = core.iram.not_i[1]
* NET 2783 = core.iram.not_aux99
* NET 2785 = core.iram.nao22_x1_3_sig
* NET 2790 = zero_to_pads
* NET 2792 = core.ialu.o3_x2_6_sig
* NET 2798 = core.ialu.na2_x1_4_sig
* NET 2799 = core.ialu.na2_x1_4_ins.i0
* NET 2800 = core.ialu.aux39
* NET 2801 = core.iram.ab_data_idx_12[3]
* NET 2802 = core.iram.ab_data_idx_9[3]
* NET 2803 = core.iram.na3_x1_60_sig
* NET 2804 = core.iram.na3_x1_61_sig
* NET 2806 = core.iram.ab_data_idx_13[3]
* NET 2809 = core.iram.aux107
* NET 2812 = core.iram.aux105
* NET 2814 = core.iram.aux112
* NET 2817 = core.iram.not_aux104
* NET 2821 = core.iram.not_aux108
* NET 2823 = core.iram.not_aux106
* NET 2825 = core.iram.aux113
* NET 2826 = core.iram.ab_data_idx_1[3]
* NET 2828 = core.iram.na3_x1_65_ins.i0
* NET 2829 = core.iram.na3_x1_64_sig
* NET 2830 = core.iram.na3_x1_63_sig
* NET 2831 = core.iram.na3_x1_62_sig
* NET 2832 = core.iram.na3_x1_65_sig
* NET 2834 = core.iram.a3_x2_14_sig
* NET 2835 = core.iram.a4_x2_4_sig
* NET 2836 = core.iram.a2_x2_14_sig
* NET 2837 = core.iram.noa2a2a2a24_x1_10_sig
* NET 2839 = core.iram.a2_x2_13_sig
* NET 2840 = core.iram.not_aux149
* NET 2841 = core.iram.not_aux128
* NET 2842 = core.iram.na2_x1_30_sig
* NET 2844 = core.iram.aux67
* NET 2846 = core.iram.ab_data_idx_6[3]
* NET 2848 = core.iram.ab_data_idx_6_3_ins.sff_s
* NET 2849 = core.iram.ab_data_idx_6_3_ins.y
* NET 2850 = core.iram.ao22_x2_28_sig
* NET 2853 = core.iram.ab_data_idx_6_3_ins.sff_m
* NET 2855 = core.iram.ab_data_idx_6_3_ins.u
* NET 2856 = core.iram.ab_data_idx_6_3_ins.ckr
* NET 2857 = core.iram.ab_data_idx_6_3_ins.nckr
* NET 2858 = p_a1.80onymous_
* NET 2859 = p_a1.57onymous_
* NET 2860 = p_np.n16c
* NET 2868 = core.ialu.aux99
* NET 2869 = core.ialu.inv_x2_9_sig
* NET 2876 = core.ialu.not_aux80
* NET 2878 = core.ialu.na2_x1_6_sig
* NET 2881 = core.ialu.not_aux33_ins.i0
* NET 2886 = core.ialu.nxr2_x1_ins.i1
* NET 2890 = core.ialu.nxr2_x1_sig
* NET 2898 = core.ialu.not_aux79
* NET 2900 = core.ialu.a2_x2_9_sig
* NET 2905 = core.ialu.o3_x2_3_sig
* NET 2907 = core.ialu.o2_x2_4_sig
* NET 2913 = core.ialu.a2_x2_7_sig
* NET 2916 = core.ialu.not_aux52
* NET 2919 = core.ialu.not_aux38
* NET 2924 = core.iram.aux111
* NET 2925 = cin_from_pads
* NET 2929 = a_from_pads[2]
* NET 2930 = a_from_pads[3]
* NET 2932 = core.iram.not_aux110
* NET 2934 = core.iram.aux115
* NET 2937 = core.iram.not_a[3]
* NET 2944 = core.ialu.xr2_x1_5_sig
* NET 2951 = core.imuxs.inv_x2_3_sig
* NET 2954 = core.imuxs.inv_x2_4_sig
* NET 2957 = core.imuxs.nao2o22_x1_2_sig
* NET 2959 = core.imuxs.y_1_ins.nq
* NET 2963 = core.imuxs.inv_x2_2_sig
* NET 2966 = core.imuxs.nao2o22_x1_sig
* NET 2968 = core.imuxs.y_0_ins.nq
* NET 2970 = core.imuxs.shift_l_ins.i0
* NET 2974 = shift_l
* NET 2975 = p_a1.1280ymous_
* NET 2976 = p_a1.cpb
* NET 2977 = p_a1.324nymous_
* NET 2979 = p_np.p6c
* NET 2980 = p_np.301nymous_
* NET 2981 = p_np.307nymous_
* NET 2982 = p_np.274nymous_
* NET 3025 = p_a1.259nymous_
* NET 3026 = p_np.997nymous_
* NET 3027 = np
* NET 3028 = p_np.cnbb
* NET 3029 = p_np.224nymous_
* NET 3030 = p_np.193nymous_
* NET 3031 = core.ialu.not_aux81_ins.i0
* NET 3034 = core.ialu.nao2o22_x1_6_sig
* NET 3038 = core.ialu.inv_x2_8_sig
* NET 3044 = core.ialu.inv_x2_7_sig
* NET 3045 = core.ialu.not_aux81
* NET 3048 = core.ialu.na2_x1_7_sig
* NET 3049 = core.ialu.na3_x1_16_ins.i0
* NET 3052 = core.ialu.na3_x1_16_sig
* NET 3053 = core.ialu.na3_x1_15_sig
* NET 3064 = core.ialu.na2_x1_5_sig
* NET 3065 = core.ialu.oa2a2a23_x2_sig
* NET 3066 = core.ialu.na3_x1_13_sig
* NET 3070 = core.ialu.not_aux39
* NET 3073 = core.ialu.aux91
* NET 3077 = core.ialu.o3_x2_2_ins.i0
* NET 3078 = core.ialu.not_aux76
* NET 3082 = core.ialu.na3_x1_6_sig
* NET 3083 = core.ialu.o3_x2_2_sig
* NET 3084 = core.ialu.alu_out_0_ins.cmd0
* NET 3085 = core.ialu.nao2o22_x1_4_sig
* NET 3098 = core.ialu.o3_x2_sig
* NET 3103 = core.ialu.not_aux1
* NET 3105 = core.ialu.o2_x2_8_sig
* NET 3106 = core.ialu.xr2_x1_4_sig
* NET 3109 = core.ialu.nxr2_x1_3_sig
* NET 3110 = core.ialu.aux3
* NET 3111 = core.rb[2]
* NET 3112 = core.imuxe.na3_x1_4_sig
* NET 3113 = core.imuxe.na2_x1_4_sig
* NET 3114 = core.imuxe.o2_x2_sig
* NET 3117 = core.imuxe.na2_x1_3_sig
* NET 3118 = core.rb[0]
* NET 3119 = core.imuxe.na3_x1_sig
* NET 3120 = core.imuxe.na2_x1_sig
* NET 3122 = core.imuxe.on12_x1_sig
* NET 3123 = core.imuxe.na3_x1_2_sig
* NET 3124 = core.imuxe.on12_x1_2_sig
* NET 3127 = core.imuxs.nao2o22_x1_3_sig
* NET 3128 = core.imuxs.y_2_ins.nq
* NET 3131 = core.imuxs.oe_ins.q
* NET 3132 = p_a1.1066ymous_
* NET 3134 = p_a1.n14c
* NET 3136 = a[1]
* NET 3137 = p_np.811nymous_
* NET 3142 = core.ialu.xr2_x1_10_sig
* NET 3144 = core.ialu.oa2a22_x2_2_ins.i3
* NET 3145 = core.ialu.xr2_x1_11_sig
* NET 3152 = core.ialu.oa2a22_x2_2_sig
* NET 3153 = core.ialu.mx3_x2_5_sig
* NET 3158 = core.ialu.oa22_x2_3_sig
* NET 3161 = core.ialu.noa22_x1_5_sig
* NET 3164 = core.ialu.no3_x1_6_sig
* NET 3165 = core.ialu.oa2ao222_x2_sig
* NET 3171 = core.ialu.aux109_ins.i0
* NET 3174 = core.ialu.na3_x1_12_sig
* NET 3177 = core.ialu.no4_x1_3_sig
* NET 3181 = core.ialu.no4_x1_sig
* NET 3188 = np_to_pads
* NET 3189 = core.ialu.na3_x1_5_sig
* NET 3194 = core.ialu.mx3_x2_sig
* NET 3200 = core.ialu.mx2_x2_sig
* NET 3209 = core.ialu.not_aux93
* NET 3218 = core.ra[2]
* NET 3220 = core.imuxe.inv_x2_2_sig
* NET 3221 = core.ra[0]
* NET 3225 = core.imuxe.inv_x2_sig
* NET 3226 = core.alu_out[0]
* NET 3230 = core.iram.r3_to_ins.q
* NET 3232 = core.iram.a2_x2_15_sig
* NET 3235 = p_ng.n18f
* NET 3239 = core.ialu.aux100
* NET 3253 = core.ialu.o3_x2_6_ins.i0
* NET 3254 = core.ialu.inv_x2_4_sig
* NET 3258 = core.ialu.o3_x2_4_sig
* NET 3260 = core.ialu.o2_x2_5_sig
* NET 3269 = core.ialu.inv_x2_5_sig
* NET 3276 = core.ialu.not_aux93_ins.i1
* NET 3277 = core.ialu.xr2_x1_3_sig
* NET 3289 = core.rb[3]
* NET 3299 = core.iram.a2_x2_15_ins.i1
* NET 3300 = p_a0.132nymous_
* NET 3301 = p_ng.n15d
* NET 3303 = core.ialu.mx3_x2_6_sig
* NET 3310 = core.ialu.aux109
* NET 3312 = core.ialu.mx2_x2_2_sig
* NET 3313 = core.ialu.inv_x2_10_sig
* NET 3319 = core.ialu.nao2o22_x1_3_sig
* NET 3322 = core.ialu.nao2o22_x1_2_sig
* NET 3325 = core.ialu.not_aux63
* NET 3327 = core.ialu.nao22_x1_8_ins.i2
* NET 3329 = core.ialu.noa22_x1_4_sig
* NET 3331 = core.ialu.aux63
* NET 3336 = core.ialu.no3_x1_7_sig
* NET 3341 = core.ialu.no4_x1_5_sig
* NET 3344 = core.ialu.o4_x2_ins.i1
* NET 3345 = core.ialu.not_aux9
* NET 3352 = core.ialu.a2_x2_8_sig
* NET 3353 = core.ialu.not_aux8
* NET 3355 = core.ialu.aux12
* NET 3362 = core.ialu.mx3_x2_3_ins.cmd1
* NET 3367 = core.ialu.aux1
* NET 3370 = core.ialu.xr2_x1_8_sig
* NET 3372 = core.ialu.xr2_x1_9_sig
* NET 3376 = core.imuxe.na3_x1_3_ins.i1
* NET 3377 = core.rb[1]
* NET 3378 = core.imuxe.na3_x1_3_sig
* NET 3379 = core.imuxe.na2_x1_2_sig
* NET 3380 = core.ra[1]
* NET 3386 = core.imuxe.a3_x2_sig
* NET 3389 = core.imuxe.not_i[2]
* NET 3390 = core.imuxs.not_noe
* NET 3391 = core.imuxs.y_3_ins.nq
* NET 3394 = core.imuxs.nao22_x1_sig
* NET 3396 = core.imuxs.inv_x2_7_sig
* NET 3397 = core.imuxs.not_aux1
* NET 3398 = core.imuxs.not_aux1_ins.i0
* NET 3399 = core.imuxs.not_aux1_ins.i1
* NET 3404 = core.imuxs.inv_x2_sig
* NET 3405 = p_a0.93onymous_
* NET 3406 = p_a0.p1
* NET 3407 = p_ng.406nymous_
* NET 3408 = p_ng.n16d
* NET 3431 = core.ialu.aux75
* NET 3445 = core.imuxe.aux3
* NET 3447 = core.imuxe.aux5
* NET 3450 = p_a0.1280ymous_
* NET 3451 = p_a0.cpb
* NET 3452 = p_a0.414nymous_
* NET 3453 = p_a0.n8b
* NET 3455 = p_ng.299nymous_
* NET 3456 = p_ng.p7a
* NET 3457 = p_ng.293nymous_
* NET 3460 = core.ialu.xr2_x1_12_sig
* NET 3468 = core.ialu.o2_x2_sig
* NET 3470 = core.ialu.a3_x2_2_sig
* NET 3477 = core.ialu.nxr2_x1_2_ins.i1
* NET 3479 = core.ialu.nxr2_x1_2_sig
* NET 3481 = core.ialu.oa22_x2_2_sig
* NET 3486 = core.ialu.a2_x2_5_sig
* NET 3488 = core.ialu.ao22_x2_4_sig
* NET 3489 = core.ialu.no3_x1_5_sig
* NET 3492 = core.ialu.aux68
* NET 3493 = ng_to_pads
* NET 3495 = core.ialu.noa22_x1_3_sig
* NET 3496 = core.ialu.na2_x1_3_sig
* NET 3499 = core.ialu.not_aux113
* NET 3502 = core.ialu.not_i_1_ins.i
* NET 3503 = core.ialu.not_aux32
* NET 3506 = core.ialu.o4_x2_sig
* NET 3507 = core.ialu.na3_x1_10_sig
* NET 3509 = core.ialu.aux4
* NET 3514 = core.ialu.not_aux5
* NET 3521 = core.ialu.not_aux89
* NET 3526 = core.ialu.not_aux67
* NET 3531 = core.ialu.a2_x2_3_sig
* NET 3532 = core.ialu.aux7
* NET 3537 = core.ialu.not_aux3
* NET 3538 = core.ialu.xr2_x1_6_sig
* NET 3548 = core.ialu.xr2_x1_7_sig
* NET 3553 = core.imuxe.not_aux0
* NET 3554 = core.imuxe.not_i[1]
* NET 3555 = core.imuxe.not_i[0]
* NET 3559 = i_from_pads[1]
* NET 3560 = core.ra[3]
* NET 3561 = core.imuxs.inv_x2_6_sig
* NET 3562 = core.imuxs.inv_x2_5_sig
* NET 3563 = core.imuxs.na4_x1_sig
* NET 3569 = core.imuxs.shift_r_ins.i0
* NET 3570 = core.imuxs.not_i[2]
* NET 3572 = p_a0.259nymous_
* NET 3573 = ng
* NET 3574 = p_ng.p3
* NET 3575 = p_ng.n5a
* NET 3576 = p_ng.n3
* NET 3577 = p_ng.224nymous_
* NET 3578 = core.ialu.not_aux101
* NET 3583 = core.ialu.not_aux74
* NET 3584 = core.ialu.aux70
* NET 3586 = core.ialu.noa3ao322_x1_ins.i6
* NET 3587 = core.ialu.inv_x2_3_sig
* NET 3591 = core.ialu.on12_x1_sig
* NET 3592 = core.ialu.not_aux68
* NET 3594 = core.ialu.not_aux56_ins.i1
* NET 3595 = core.ialu.no2_x1_6_sig
* NET 3599 = core.ialu.not_aux56
* NET 3602 = core.ialu.nao22_x1_8_sig
* NET 3603 = core.ialu.na3_x1_9_sig
* NET 3604 = core.ialu.nao22_x1_7_sig
* NET 3606 = core.ialu.no4_x1_2_sig
* NET 3608 = core.ialu.no2_x1_5_sig
* NET 3611 = core.ialu.na3_x1_8_sig
* NET 3613 = core.ialu.noa22_x1_sig
* NET 3614 = core.ialu.not_aux15
* NET 3616 = core.ialu.no2_x1_2_sig
* NET 3619 = core.ialu.not_aux0
* NET 3621 = core.ialu.no2_x1_sig
* NET 3622 = core.ialu.na3_x1_11_sig
* NET 3623 = core.ialu.not_aux13
* NET 3624 = core.ialu.na3_x1_4_sig
* NET 3625 = core.ialu.na3_x1_3_sig
* NET 3627 = core.ialu.a3_x2_3_ins.i0
* NET 3629 = core.ialu.a3_x2_3_sig
* NET 3630 = core.ialu.nao22_x1_6_sig
* NET 3634 = core.ialu.no2_x1_7_sig
* NET 3635 = core.s[0]
* NET 3636 = core.ialu.not_r[0]
* NET 3637 = core.ialu.not_s[0]
* NET 3638 = core.r[0]
* NET 3639 = core.imuxe.na3_x1_5_sig
* NET 3641 = core.imuxe.on12_x1_4_sig
* NET 3642 = core.imuxe.on12_x1_3_sig
* NET 3643 = core.imuxe.not_aux1
* NET 3645 = core.imuxe.na2_x1_5_sig
* NET 3646 = core.imuxe.not_aux4
* NET 3647 = i_from_pads[2]
* NET 3650 = core.imuxe.aux2
* NET 3651 = core.imuxe.inv_x2_3_sig
* NET 3655 = core.saccu[0]
* NET 3659 = core.iaccu.na2_x1_4_ins.i0
* NET 3660 = p_a0.196nymous_
* NET 3661 = a_from_pads[0]
* NET 3662 = a[0]
* NET 3663 = p_ng.889nymous_
* NET 3664 = p_ng.793nymous_
* NET 3686 = p_a0.n14a
* NET 3687 = p_a0.568nymous_
* NET 3690 = core.ialu.not_aux107_ins.i0
* NET 3691 = core.ialu.a2_x2_11_sig
* NET 3694 = core.ialu.not_aux107
* NET 3700 = core.ialu.noa3ao322_x1_sig
* NET 3701 = core.ialu.nao22_x1_5_sig
* NET 3710 = core.r[3]
* NET 3712 = core.s[3]
* NET 3714 = core.ialu.aux42
* NET 3715 = ovr_to_pads
* NET 3716 = core.ialu.na3_x1_2_sig
* NET 3717 = core.ialu.ovr_ins.i0
* NET 3724 = core.ialu.na4_x1_sig
* NET 3726 = core.ialu.nao22_x1_3_sig
* NET 3727 = core.ialu.aux16
* NET 3729 = core.ialu.ao22_x2_sig
* NET 3732 = core.ialu.nao22_x1_sig
* NET 3733 = core.ialu.ao2o22_x2_sig
* NET 3740 = core.ialu.na3_x1_7_sig
* NET 3742 = core.ialu.o2_x2_2_sig
* NET 3744 = core.ialu.a2_x2_6_sig
* NET 3748 = core.ialu.mx3_x2_3_sig
* NET 3760 = core.ialu.a4_x2_sig
* NET 3766 = core.ialu.na3_x1_sig
* NET 3771 = core.ialu.na2_x1_sig
* NET 3772 = core.ialu.na2_x1_2_sig
* NET 3774 = core.ialu.not_aux78
* NET 3781 = core.ialu.not_aux37
* NET 3785 = core.ialu.a2_x2_sig
* NET 3786 = core.ialu.not_aux7
* NET 3792 = core.saccu[3]
* NET 3793 = core.imuxe.not_accu[2]
* NET 3797 = core.iaccu.a2_x2_sig
* NET 3798 = core.iaccu.a2_x2_ins.i0
* NET 3799 = core.imuxe.inv_x2_4_sig
* NET 3804 = core.iaccu.no2_x1_5_sig
* NET 3806 = core.iaccu.nao22_x1_2_sig
* NET 3813 = core.iaccu.na2_x1_4_sig
* NET 3814 = core.iaccu.oa22_x2_4_sig
* NET 3819 = core.ialu.o3_x2_11_ins.i1
* NET 3823 = core.ialu.o3_x2_7_sig
* NET 3824 = core.ialu.oa22_x2_4_sig
* NET 3825 = core.ialu.o2_x2_9_sig
* NET 3829 = core.ialu.aux32
* NET 3832 = core.ialu.o2_x2_10_sig
* NET 3833 = core.ialu.na3_x1_17_sig
* NET 3835 = core.alu_out[3]
* NET 3839 = core.ialu.not_aux33
* NET 3840 = core.ialu.not_aux41
* NET 3843 = core.ialu.no3_x1_2_sig
* NET 3844 = core.ialu.nao22_x1_2_sig
* NET 3846 = core.ialu.not_i[1]
* NET 3847 = core.ialu.noa22_x1_2_sig
* NET 3851 = core.ialu.no2_x1_8_sig
* NET 3852 = core.ialu.ao22_x2_2_sig
* NET 3855 = core.ialu.na3_x1_14_sig
* NET 3858 = core.ialu.o2_x2_6_sig
* NET 3861 = core.ialu.o2_x2_7_sig
* NET 3864 = core.ialu.o2_x2_3_sig
* NET 3865 = core.ialu.ao2o22_x2_2_sig
* NET 3871 = core.ialu.not_aux110
* NET 3872 = core.ialu.mx3_x2_4_sig
* NET 3880 = core.ialu.inv_x2_6_sig
* NET 3881 = core.ialu.oa2a22_x2_sig
* NET 3882 = core.ialu.not_aux4
* NET 3884 = core.ialu.oa2a22_x2_ins.i0
* NET 3886 = core.ialu.not_aux77
* NET 3887 = core.ialu.mx3_x2_2_sig
* NET 3895 = core.ialu.nao2o22_x1_5_ins.i3
* NET 3896 = core.ialu.nao2o22_x1_5_sig
* NET 3902 = core.ialu.aux98
* NET 3904 = core.saccu[2]
* NET 3905 = core.alu_out[1]
* NET 3907 = core.saccu[1]
* NET 3908 = core.iaccu.no2_x1_3_ins.i0
* NET 3911 = core.alu_out[2]
* NET 3914 = core.iaccu.not_aux4_ins.i1
* NET 3916 = core.iaccu.not_i[2]
* NET 3917 = core.iaccu.inv_x2_2_sig
* NET 3918 = core.iaccu.accu_reg[3]
* NET 3920 = core.iaccu.accu_reg_3_ins.sff_s
* NET 3921 = core.iaccu.na3_x1_4_sig
* NET 3922 = core.iaccu.accu_reg_3_ins.y
* NET 3925 = core.iaccu.accu_reg_3_ins.sff_m
* NET 3926 = core.iaccu.accu_reg_3_ins.ck
* NET 3927 = core.iaccu.accu_reg_3_ins.u
* NET 3928 = core.iaccu.accu_reg_3_ins.nckr
* NET 3929 = core.iaccu.accu_reg_3_ins.ckr
* NET 3930 = p_q0.eb
* NET 3931 = q0_to_pads
* NET 3932 = p_q0.126nymous_
* NET 3933 = p_q3.n17d
* NET 3968 = p_q0.50onymous_
* NET 3969 = p_q0.472nymous_
* NET 3970 = p_q3.n16d
* NET 3971 = p_q3.32onymous_
* NET 3972 = core.ialu.nao22_x1_9_sig
* NET 3973 = core.ialu.o3_x2_11_sig
* NET 3977 = core.ialu.a2_x2_10_sig
* NET 3980 = core.ialu.an12_x1_sig
* NET 3981 = core.ialu.oa2a2a2a24_x2_sig
* NET 3982 = core.ialu.na2_x1_10_sig
* NET 3983 = core.ialu.not_s[2]
* NET 3986 = core.ialu.o3_x2_9_sig
* NET 3990 = core.ialu.o2_x2_11_ins.i1
* NET 3991 = core.s[2]
* NET 3993 = core.ialu.o2_x2_11_sig
* NET 3994 = core.ialu.not_aux43
* NET 3996 = core.ialu.oa22_x2_sig
* NET 4001 = core.ialu.no2_x1_3_sig
* NET 4003 = core.ialu.inv_x2_11_sig
* NET 4005 = core.ialu.not_aux112
* NET 4008 = core.ialu.not_aux115
* NET 4010 = core.ialu.not_aux49
* NET 4016 = core.ialu.aux77
* NET 4020 = core.ialu.a2_x2_4_sig
* NET 4024 = core.ialu.not_aux47
* NET 4028 = core.ialu.a2_x2_2_sig
* NET 4032 = core.ialu.aux19
* NET 4034 = core.ialu.not_aux95
* NET 4039 = core.ialu.not_s[1]
* NET 4044 = core.iaccu.na2_x1_2_sig
* NET 4051 = core.iaccu.oa22_x2_2_sig
* NET 4053 = core.iaccu.no2_x1_2_sig
* NET 4054 = core.iaccu.o3_x2_2_sig
* NET 4056 = core.iaccu.no2_x1_3_sig
* NET 4058 = core.iaccu.not_aux4
* NET 4059 = core.iaccu.no2_x1_sig
* NET 4065 = core.iaccu.o2_x2_sig
* NET 4067 = core.iaccu.not_aux0
* NET 4068 = core.iaccu.o3_x2_4_sig
* NET 4071 = q3_from_pads
* NET 4072 = core.iaccu.no2_x1_4_sig
* NET 4075 = p_q0.n6a
* NET 4076 = p_q0.1292ymous_
* NET 4077 = p_q0.329nymous_
* NET 4078 = p_q0.330nymous_
* NET 4079 = p_q3.p6a
* NET 4080 = p_q3.57onymous_
* NET 4081 = p_q3.53onymous_
* NET 4082 = p_q3.113nymous_
* NET 4083 = p_q3.n0
* NET 4084 = q3_to_pads
* NET 4090 = core.ialu.not_aux103
* NET 4092 = core.ialu.na2_x1_11_sig
* NET 4094 = core.ialu.inv_x2_12_sig
* NET 4096 = core.ialu.aux102
* NET 4098 = core.ialu.aux51
* NET 4101 = core.ialu.a3_x2_ins.i0
* NET 4102 = core.ialu.ao22_x2_3_ins.i2
* NET 4104 = core.ialu.aux105
* NET 4105 = core.ialu.not_cin
* NET 4107 = core.ialu.o3_x2_5_ins.i2
* NET 4111 = core.ialu.on12_x1_2_sig
* NET 4117 = core.iaccu.not_aux2_ins.i0
* NET 4118 = core.iaccu.accu_reg_0_ins.ck
* NET 4119 = core.iaccu.na2_x1_ins.i0
* NET 4121 = p_q3.612nymous_
* NET 4122 = core.iaccu.o3_x2_sig
* NET 4123 = core.iaccu.na2_x1_sig
* NET 4124 = p_q0.265nymous_
* NET 4125 = q0
* NET 4126 = p_q3.784nymous_
* NET 4127 = p_q3.898nymous_
* NET 4128 = q3
* NET 4129 = p_q3.162nymous_
* NET 4130 = p_q3.778nymous_
* NET 4132 = core.ialu.o3_x2_10_sig
* NET 4135 = core.ialu.o3_x2_12_sig
* NET 4137 = core.ialu.not_aux40
* NET 4139 = core.ialu.no2_x1_9_sig
* NET 4142 = core.ialu.a3_x2_sig
* NET 4143 = core.ialu.aux43_ins.i0
* NET 4144 = core.ialu.aux43
* NET 4146 = core.ialu.not_aux60
* NET 4148 = core.ialu.not_aux62
* NET 4150 = core.ialu.nao22_x1_4_sig
* NET 4152 = core.ialu.ao22_x2_3_sig
* NET 4157 = core.ialu.no3_x1_4_sig
* NET 4161 = core.ialu.not_aux106
* NET 4163 = core.ialu.not_aux42
* NET 4164 = core.ialu.nao2o22_x1_sig
* NET 4167 = core.ialu.not_aux105
* NET 4169 = core.ialu.no4_x1_4_sig
* NET 4174 = core.ialu.o3_x2_5_sig
* NET 4177 = core.ialu.not_aux28
* NET 4179 = core.ialu.aux29
* NET 4182 = core.ialu.not_aux31
* NET 4186 = core.ialu.not_aux54
* NET 4187 = core.ialu.not_r[1]
* NET 4191 = core.ialu.xr2_x1_2_sig
* NET 4196 = core.s[1]
* NET 4198 = core.r[1]
* NET 4202 = core.iaccu.accu_reg_1_ins.ckr
* NET 4203 = core.iaccu.accu_reg_1_ins.nckr
* NET 4205 = core.iaccu.accu_reg_1_ins.sff_s
* NET 4206 = core.iaccu.accu_reg_1_ins.sff_m
* NET 4208 = core.iaccu.accu_reg_1_ins.y
* NET 4210 = core.iaccu.na3_x1_2_sig
* NET 4211 = core.iaccu.accu_reg_1_ins.u
* NET 4213 = core.iaccu.not_aux2
* NET 4214 = core.iaccu.accu_reg[0]
* NET 4215 = core.iaccu.accu_reg_0_ins.ckr
* NET 4216 = core.iaccu.accu_reg_0_ins.nckr
* NET 4217 = core.iaccu.accu_reg_0_ins.sff_m
* NET 4219 = core.iaccu.accu_reg_0_ins.y
* NET 4220 = core.iaccu.accu_reg_0_ins.sff_s
* NET 4221 = core.iaccu.na3_x1_sig
* NET 4224 = core.iaccu.accu_reg_0_ins.u
* NET 4229 = p_q0.nt
* NET 4230 = p_q0.n14b
* NET 4231 = p_q0.208nymous_
* NET 4233 = core.ialu.not_aux50
* NET 4236 = core.ialu.o2_x2_13_sig
* NET 4238 = core.ialu.na3_x1_20_sig
* NET 4240 = core.ialu.not_aux104
* NET 4241 = core.ialu.aux104
* NET 4243 = core.ialu.not_i[0]
* NET 4246 = core.ialu.a2_x2_12_sig
* NET 4247 = core.ialu.na2_x1_9_sig
* NET 4248 = core.ialu.na2_x1_8_sig
* NET 4250 = core.ialu.na3_x1_18_sig
* NET 4253 = core.ialu.aux108_ins.i0
* NET 4256 = core.ialu.na4_x1_2_sig
* NET 4258 = core.ialu.aux108
* NET 4259 = core.ialu.aux114
* NET 4260 = core.ialu.inv_x2_2_sig
* NET 4261 = core.ialu.not_aux102
* NET 4263 = core.ialu.no2_x1_4_sig
* NET 4264 = core.ialu.no3_x1_3_sig
* NET 4265 = core.ialu.na3_x1_19_sig
* NET 4266 = core.ialu.o3_x2_8_sig
* NET 4269 = core.ialu.not_i[2]
* NET 4270 = core.ialu.o2_x2_12_sig
* NET 4272 = core.ialu.not_aux61
* NET 4273 = core.ialu.not_aux17
* NET 4275 = core.ialu.na4_x1_3_sig
* NET 4278 = core.ialu.aux111
* NET 4279 = core.ialu.not_aux69
* NET 4280 = core.ialu.not_aux48
* NET 4283 = core.ialu.not_aux16
* NET 4284 = core.ialu.aux17
* NET 4285 = core.ialu.not_aux21
* NET 4287 = core.ialu.not_aux19
* NET 4289 = core.ialu.aux21
* NET 4290 = core.ialu.aux25_ins.i0
* NET 4292 = core.ialu.aux25
* NET 4293 = core.ialu.inv_x2_sig
* NET 4295 = core.ialu.not_aux22
* NET 4296 = core.ialu.no3_x1_sig
* NET 4297 = core.ialu.not_aux24
* NET 4298 = core.ialu.aux23
* NET 4301 = core.ialu.aux20
* NET 4302 = core.ialu.not_aux20
* NET 4303 = core.ialu.not_aux23
* NET 4305 = core.ialu.not_aux97
* NET 4308 = core.ialu.xr2_x1_sig
* NET 4311 = core.iaccu.accu_reg_2_ins.sff_s
* NET 4312 = core.iaccu.accu_reg_2_ins.y
* NET 4313 = core.iaccu.accu_reg_2_ins.sff_m
* NET 4317 = core.iaccu.accu_reg_2_ins.nckr
* NET 4318 = core.iaccu.accu_reg_2_ins.u
* NET 4319 = core.iaccu.accu_reg_2_ins.ckr
* NET 4320 = core.iaccu.not_accu_reg[2]
* NET 4322 = core.iaccu.accu_reg[2]
* NET 4324 = core.iaccu.o3_x2_3_sig
* NET 4325 = core.iaccu.na2_x1_3_sig
* NET 4327 = core.iaccu.na3_x1_3_sig
* NET 4329 = core.iaccu.accu_reg[1]
* NET 4332 = core.iaccu.oa22_x2_3_sig
* NET 4334 = core.iaccu.not_accu_reg[3]
* NET 4337 = core.iaccu.not_aux3
* NET 4338 = core.iaccu.not_aux1
* NET 4339 = core.iaccu.o2_x2_2_sig
* NET 4341 = core.iaccu.inv_x2_sig
* NET 4342 = q0_from_pads
* NET 4343 = core.iaccu.oa22_x2_sig
* NET 4345 = core.iaccu.not_i[1]
* NET 4346 = core.iaccu.nao22_x1_sig
* NET 4347 = core.iaccu.not_accu_reg[1]
* NET 4350 = r3_from_pads
* NET 4352 = shift_r
* NET 4354 = p_r0.126nymous_
* NET 4355 = p_r3.n17d
* NET 4356 = p_r0.538nymous_
* NET 4357 = p_r0.64onymous_
* NET 4358 = p_r3.n16c
* NET 4359 = p_r3.25onymous_
* NET 4360 = p_r0.1292ymous_
* NET 4361 = p_r0.cpb
* NET 4362 = p_r0.329nymous_
* NET 4363 = p_r0.330nymous_
* NET 4364 = p_r3.p6a
* NET 4365 = p_r3.57onymous_
* NET 4366 = p_r3.53onymous_
* NET 4367 = p_r3.n2
* NET 4369 = p_r0.265nymous_
* NET 4370 = p_r3.784nymous_
* NET 4371 = r3
* NET 4373 = p_r3.cnbb
* NET 4376 = p_r0.1078ymous_
* NET 4378 = p_r0.n14b
* NET 4380 = r0
* NET 4381 = p_r3.914nymous_
* NET 4382 = p_cout.n18d
* NET 4383 = p_cin.p0
* NET 4384 = p_cout.n15d
* NET 4385 = p_cin.n1
* NET 4386 = p_cin.p1
* NET 4387 = p_cin.p12
* NET 4388 = p_cout.406nymous_
* NET 4389 = p_cout.n16d
* NET 4390 = p_cin.1280ymous_
* NET 4391 = p_cin.cpb
* NET 4392 = p_cin.n8b
* NET 4394 = p_cout.299nymous_
* NET 4395 = p_cout.p7a
* NET 4396 = p_cout.293nymous_
* NET 4397 = cout_to_pads
* NET 4398 = p_cin.259nymous_
* NET 4399 = p_cout.227nymous_
* NET 4400 = cout
* NET 4401 = p_cout.p3
* NET 4402 = p_cout.n5a
* NET 4403 = p_cout.n3
* NET 4404 = p_cout.224nymous_
* NET 4406 = p_cin.221nymous_
* NET 4408 = cin
* NET 4409 = p_cout.168nymous_
* NET 4410 = p_cin.n14a
* NET 4411 = p_cin.568nymous_
* NET 4413 = p_y3.144nymous_
* NET 4414 = p_y3.119nymous_
* NET 4417 = p_y3.nnt
* NET 4418 = p_y3.1062ymous_
* NET 4420 = p_y2.p3
* NET 4421 = p_y2.131nymous_
* NET 4425 = p_y2.257nymous_
* NET 4426 = p_y2.219nymous_
* NET 4428 = p_y1.111nymous_
* NET 4430 = p_y1.99onymous_
* NET 4431 = p_y1.638nymous_
* NET 4432 = p_y1.43onymous_
* NET 4433 = p_y1.257nymous_
* NET 4434 = p_y1.nt
* NET 4435 = p_y1.969nymous_
* NET 4438 = p_y0.119nymous_
* NET 4440 = p_y0.80onymous_
* NET 4441 = p_y0.257nymous_
* NET 4442 = p_y0.1062ymous_
* NET 4444 = p_vssick0.230nymous_
* NET 4445 = p_vsseck1.31onymous_
* NET 4446 = p_vsseck0.31onymous_
* NET 4447 = p_d3.p3
* NET 4448 = p_d3.132nymous_
* NET 4449 = p_d3.p1
* NET 4450 = p_d3.259nymous_
* NET 4451 = p_d3.196nymous_
* NET 4452 = d_from_pads[3]
* NET 4453 = p_d2.112nymous_
* NET 4454 = p_d2.640nymous_
* NET 4455 = p_d2.43onymous_
* NET 4456 = p_d2.nnt
* NET 4457 = p_d2.nt
* NET 4458 = d_from_pads[2]
* NET 4459 = p_d1.639nymous_
* NET 4460 = p_d1.132nymous_
* NET 4461 = p_d1.532nymous_
* NET 4462 = p_d1.259nymous_
* NET 4463 = p_d1.1066ymous_
* NET 4464 = d_from_pads[1]
* NET 4465 = p_d0.639nymous_
* NET 4466 = p_d0.p0
* NET 4467 = p_d0.p1
* NET 4468 = p_d0.259nymous_
* NET 4469 = p_d0.221nymous_
* NET 4470 = d_from_pads[0]
* NET 4476 = ck_ring
* NET 4478 = vddi
* NET 4479 = p_y3.1275ymous_
* NET 4480 = p_y3.cpb
* NET 4481 = p_y2.cpb
* NET 4482 = p_y2.1275ymous_
* NET 4483 = p_y1.n6a
* NET 4484 = p_y1.1275ymous_
* NET 4485 = p_y0.1275ymous_
* NET 4486 = p_y0.cpb
* NET 4487 = p_d3.1280ymous_
* NET 4488 = p_d3.cpb
* NET 4489 = p_d2.n6a
* NET 4490 = p_d2.1280ymous_
* NET 4491 = p_d1.1280ymous_
* NET 4492 = p_d1.cpb
* NET 4493 = p_d0.1280ymous_
* NET 4494 = p_d0.cpb
* NET 4495 = p_y3.57onymous_
* NET 4496 = p_y3.1335ymous_
* NET 4498 = p_y3.n14c
* NET 4500 = p_y2.410nymous_
* NET 4501 = p_y2.1336ymous_
* NET 4503 = p_y2.n14a
* NET 4504 = p_y2.564nymous_
* NET 4505 = p_y1.459nymous_
* NET 4506 = p_y1.n8a
* NET 4507 = p_y1.319nymous_
* NET 4508 = p_y1.n14b
* NET 4509 = p_y1.201nymous_
* NET 4510 = p_y0.57onymous_
* NET 4511 = p_y0.1335ymous_
* NET 4513 = p_y0.n14c
* NET 4515 = p_d3.414nymous_
* NET 4516 = p_d3.n8b
* NET 4518 = p_d3.n14a
* NET 4519 = p_d3.568nymous_
* NET 4520 = p_d2.466nymous_
* NET 4521 = p_d2.n8a
* NET 4522 = p_d2.324nymous_
* NET 4523 = p_d2.n14b
* NET 4524 = p_d2.87onymous_
* NET 4525 = p_d1.57onymous_
* NET 4526 = p_d1.1341ymous_
* NET 4528 = p_d1.n14c
* NET 4530 = p_d0.p12
* NET 4531 = p_d0.n8b
* NET 4533 = p_d0.n14a
* NET 4534 = p_d0.568nymous_
* NET 4535 = vdde
* NET 4536 = y[3]
* NET 4537 = y[2]
* NET 4538 = y[1]
* NET 4539 = y[0]
* NET 4540 = vssi
* NET 4541 = vsse
* NET 4542 = d[3]
* NET 4543 = d[2]
* NET 4544 = d[1]
* NET 4545 = d[0]
Mtr_10362 4478 2596 2594 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10361 2495 2593 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10360 2594 2785 2495 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10359 4478 1591 1004 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10358 1004 830 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10357 4478 829 1004 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10356 1004 1564 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10355 211 365 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_10354 1972 1842 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10353 1411 1492 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_10352 825 829 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_10351 1708 1878 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10350 846 877 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10349 381 708 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_10348 2426 2802 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_10347 2092 2079 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10346 2079 2196 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10345 4478 2076 2079 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10344 2079 2075 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10343 4478 2084 2079 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10342 745 744 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10341 4478 2782 744 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10340 744 692 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10339 1119 1564 1122 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10338 1120 1118 1119 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10337 1121 1975 1120 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10336 4478 1412 1121 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10335 4478 1122 1123 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10334 2593 2590 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10333 4478 2600 2590 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10332 2590 2783 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10331 1489 1487 2111 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10330 4478 1488 1489 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10329 1697 1696 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10328 4478 3905 1697 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10327 1527 1514 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10326 4478 1516 1514 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10325 1514 1446 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10324 1552 1490 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10323 4478 2284 1490 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10322 1490 1405 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10321 328 302 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10320 4478 303 302 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10319 302 300 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10318 1706 1705 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10317 4478 2778 1706 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10316 402 403 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10315 4478 404 403 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10314 403 401 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10313 1317 1318 1321 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_10312 4478 1315 1317 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_10311 1426 1321 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10310 2620 1428 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10309 1710 1568 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10308 4478 1591 1568 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10307 1568 1569 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10306 2004 1714 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10305 4478 1710 1714 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10304 1714 1713 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10303 1730 1573 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10302 4478 1782 1573 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10301 1573 1710 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10300 4478 1492 1412 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10299 1409 1972 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10298 1412 3226 1409 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10297 4478 2929 2821 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10296 2821 2820 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10295 4478 3661 2820 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10294 2932 2929 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10293 4478 3661 2932 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10292 2410 2814 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10291 2414 2825 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_10290 1646 2934 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_10289 2816 3661 2818 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10288 4478 2929 2816 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10287 2817 2818 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10286 4478 1551 1555 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10285 1555 1556 1554 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10284 1554 1552 1553 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10283 1976 1553 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10282 404 263 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10281 4478 1591 263 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10280 263 265 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10279 238 220 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10278 4478 1564 220 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10277 220 1302 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10276 605 583 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10275 4478 581 583 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10274 583 580 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10273 1569 1566 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10272 4478 1564 1566 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10271 1566 1565 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10270 2542 2447 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10269 4478 2289 2424 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10268 2289 2285 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10267 4478 2584 2246 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10266 2246 2287 2289 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10265 4478 1834 1843 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10264 1843 1833 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10263 1843 1842 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10262 743 741 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10261 4478 689 741 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10260 741 694 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10259 510 206 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10258 4478 365 206 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10257 206 207 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10256 4478 1110 1114 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10255 1113 1835 1112 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10254 1112 1118 1116 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10253 1114 1111 1113 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10252 456 803 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10251 4478 456 457 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10250 457 459 730 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10249 4478 1782 182 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10248 183 212 479 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10247 182 211 183 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10246 1758 1754 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10245 4478 1758 1679 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10244 1679 1755 2635 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10243 2813 2817 2812 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10242 4478 2930 2813 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10241 2810 2821 2811 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10240 4478 2930 2810 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10239 2922 2932 2924 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10238 4478 2930 2922 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10237 2822 2821 2827 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10236 4478 2937 2822 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10235 2782 2766 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_10234 4478 1491 1565 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10233 1406 1407 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10232 1406 1697 1491 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10231 1491 1405 1406 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10230 1516 1493 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10229 4478 1565 1493 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10228 1493 1413 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10227 2138 2137 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10226 4478 2136 2137 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10225 2137 2139 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10224 1295 2136 1296 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_10223 4478 1301 1295 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_10222 1294 1296 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10221 406 382 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10220 4478 1294 382 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10219 382 383 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10218 633 408 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10217 4478 406 408 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10216 408 407 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10215 441 439 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10214 4478 633 439 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10213 439 438 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10212 4478 1285 1287 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10211 1285 1288 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10210 4478 1552 1286 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10209 1286 1284 1285 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10208 265 216 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10207 4478 1302 216 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10206 216 213 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10205 303 267 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10204 4478 265 267 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10203 267 264 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10202 2335 2812 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10201 4478 3661 2823 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10200 2823 2819 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10199 4478 2929 2819 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10198 2337 2809 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10197 385 235 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10196 4478 1591 235 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10195 235 406 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10194 1589 1501 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10193 4478 1591 1501 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10192 1501 1516 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10191 658 423 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10190 4478 1782 423 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10189 423 605 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10188 1804 1788 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10187 4478 1782 1788 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10186 1788 1785 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10185 2222 1911 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_10184 2220 2696 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10183 296 290 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10182 4478 291 290 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10181 290 300 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10180 581 545 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10179 4478 1564 545 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10178 545 1294 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10177 2290 1974 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10176 4478 1972 1974 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10175 1974 2778 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10174 2695 2781 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10173 4478 2323 2250 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10172 2251 2620 2301 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10171 2250 2781 2251 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10170 2529 2527 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10169 4478 2445 2527 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10168 2527 2449 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10167 898 899 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10166 4478 896 899 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10165 899 900 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10164 1921 2542 1920 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10163 4478 1919 1921 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10162 1963 2220 2094 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10161 4478 2091 1963 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10160 1912 2390 1914 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10159 4478 1913 1912 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10158 1924 2222 1923 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10157 4478 1922 1924 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10156 4478 1837 1840 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10155 1841 1838 1977 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10154 1840 2584 1841 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10153 4478 1412 694 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10152 694 1564 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10151 694 693 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10150 4478 693 692 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10149 692 1552 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10148 692 1564 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10147 4478 1150 1133 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10146 1133 1299 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10145 1133 1123 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10144 4478 1298 1150 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10143 1149 1148 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10142 1150 2171 1149 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10141 4478 1297 1299 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10140 1300 1301 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10139 1299 1298 1300 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10138 4478 1564 1293 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10137 1292 1838 1297 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10136 1293 1552 1292 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10135 4478 2582 2761 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10134 2478 2483 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10133 2761 2476 2478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10132 4478 2471 2475 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10131 2474 2806 2479 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10130 2475 2472 2474 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10129 2247 2782 2292 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10128 4478 2290 2247 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10127 2476 2292 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10126 2484 2589 2588 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10125 4478 2806 2484 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10124 2587 2588 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10123 2480 2584 2586 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10122 4478 2585 2480 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10121 2470 2778 2577 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10120 4478 2468 2470 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10119 4478 2782 2785 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10118 2784 2783 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10117 2785 3835 2784 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10116 4478 2601 2596 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10115 2596 2592 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10114 2596 2598 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10113 4478 2600 2601 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10112 2496 2620 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10111 2601 2621 2496 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10110 4478 1499 2143 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10109 2143 1564 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10108 2143 1591 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10107 999 2620 998 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10106 4478 997 999 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10105 1000 998 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10104 4478 1972 1008 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10103 1008 1009 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10102 4478 1032 1009 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10101 1006 1004 1007 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10100 4478 1552 1006 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10099 1492 2136 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10098 4478 1972 1492 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10097 2780 2778 2781 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10096 4478 2779 2780 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10095 4478 1407 1291 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_10094 1291 2782 1289 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_10093 1289 1411 1290 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_10092 1288 1290 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10091 4478 1700 1701 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10090 1702 1701 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10089 4478 1705 1701 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10088 1701 3905 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10087 4478 2284 2245 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_10086 2245 2290 2244 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_10085 2244 2782 2286 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_10084 2285 2286 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10083 786 1782 2197 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10082 4478 785 786 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10081 4478 1843 1847 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10080 1845 2138 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10079 1847 1844 1845 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10078 4478 1625 1624 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10077 1625 1627 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10076 4478 2217 1626 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10075 1626 2070 1625 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10074 4478 436 435 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10073 436 440 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10072 4478 2217 437 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10071 437 913 436 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10070 4478 325 320 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10069 325 326 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10068 4478 2217 195 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10067 195 723 325 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10066 4478 2218 2215 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10065 2218 2399 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10064 4478 2217 2219 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10063 2219 2688 2218 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10062 4478 763 543 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10061 843 543 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10060 4478 544 543 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10059 543 541 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10058 4478 855 227 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10057 375 227 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10056 4478 229 227 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10055 227 224 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10054 4478 2323 2256 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10053 2257 2325 2322 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10052 2256 2781 2257 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10051 1067 918 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10050 4478 917 918 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10049 918 1096 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10048 2087 1803 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_10047 4478 1798 1803 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10046 1803 1815 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10045 1798 1769 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10044 4478 1765 1769 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10043 1769 1764 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10042 4478 2513 1142 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10041 1142 1143 1141 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10040 1141 2423 1144 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10039 1180 1144 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10038 4478 877 887 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10037 887 1428 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10036 887 880 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10035 4478 913 888 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10034 888 2197 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10033 888 722 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10032 4478 1812 1809 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10031 1809 2696 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10030 1809 1806 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_10029 4478 1885 1789 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10028 1789 2357 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10027 1789 1774 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10026 4478 1810 1797 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10025 1797 1911 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10024 1797 1794 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10023 4478 1886 1790 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10022 1790 2656 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10021 1790 1774 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10020 1957 2325 2026 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10019 4478 2022 1957 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10018 4478 2513 1953 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10017 1953 2160 1952 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10016 1952 2423 2011 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10015 2041 2011 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_10014 4478 2070 2064 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10013 2064 2197 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10012 2064 2059 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10011 4478 1878 2035 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10010 2035 2437 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10009 2035 1879 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10008 4478 2195 2179 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10007 2179 2447 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10006 2179 2178 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10005 4478 2295 2130 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10004 2130 1985 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10003 2130 1984 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_10002 4478 1975 1944 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10001 1944 2290 1945 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_10000 1945 1976 1980 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09999 1984 1980 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09998 4478 1977 1985 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09997 1946 1981 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09996 1985 2516 1946 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09995 4478 521 516 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09994 478 515 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09993 516 2325 478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09992 1836 1835 1839 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_09991 4478 1976 1836 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_09990 2472 1839 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09989 4478 2581 2477 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09988 2582 2587 2477 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09987 2477 2586 2582 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09986 2581 2579 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09985 2473 2576 2469 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09984 2473 2577 4478 4478 tp L=0.32U W=4.05U AS=3.0375P AD=3.0375P PS=9.6U PD=9.6U 
Mtr_09983 4478 2806 2473 4478 tp L=0.32U W=4.05U AS=3.0375P AD=3.0375P PS=9.6U PD=9.6U 
Mtr_09982 2469 2620 2579 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09981 2579 2806 2473 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09980 4478 2143 2145 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09979 2145 2146 2144 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09978 2144 2147 2148 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09977 2592 2148 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09976 1013 1002 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09975 4478 1032 1003 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09974 1003 1000 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09973 1003 1116 1005 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09972 1005 1001 1003 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09971 1002 1007 1005 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09970 1005 1008 1002 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09969 1627 1896 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09968 4478 1894 1627 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09967 440 441 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09966 4478 763 440 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09965 326 328 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09964 4478 855 326 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09963 2399 2699 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09962 4478 2457 2399 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09961 2191 1895 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09960 4478 1894 2191 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09959 4478 843 762 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09958 845 846 762 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09957 762 2297 845 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09956 4478 375 379 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09955 380 381 379 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09954 379 2297 380 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09953 4478 2301 2249 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09952 2774 2426 2249 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09951 2249 2297 2774 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09950 1747 1885 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_09949 696 1051 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_09948 4478 2322 2255 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09947 2317 2320 2255 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09946 2255 2315 2317 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09945 1193 1197 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09944 4478 1192 1197 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09943 1197 1235 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09942 1192 1178 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09941 4478 1176 1178 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09940 1178 1175 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09939 917 873 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09938 4478 874 873 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09937 873 871 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09936 4478 1090 1066 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09935 1066 1911 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09934 1066 1072 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09933 4478 904 900 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09932 900 2447 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09931 900 903 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09930 4478 1160 896 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09929 896 2435 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09928 896 714 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09927 4478 1061 1062 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09926 1062 2656 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09925 1062 1072 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09924 4478 1789 2202 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09923 2202 1797 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09922 4478 1790 2202 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09921 2202 1809 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09920 4478 2041 2203 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09919 2203 2042 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09918 4478 2043 2203 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09917 2203 2044 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09916 1961 2513 2031 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09915 4478 2032 1961 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09914 4478 2516 2295 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09913 2248 2307 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09912 2295 2325 2248 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09911 2008 2055 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_09910 603 614 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09909 4478 763 603 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09908 288 296 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09907 4478 855 288 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09906 2366 2699 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09905 4478 2544 2366 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09904 1642 1472 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09903 4478 1894 1642 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09902 859 1347 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09901 2320 2356 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_09900 1846 1849 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09899 4478 1846 1848 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09898 1848 1847 1894 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09897 763 761 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09896 4478 1287 761 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09895 761 698 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09894 1304 2284 1303 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09893 4478 1301 1304 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09892 1302 1303 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09891 4478 1702 1667 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09890 1704 1706 1667 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09889 1667 2782 1704 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09888 855 849 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09887 4478 1704 849 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09886 849 848 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09885 2514 2781 2617 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09884 4478 2513 2514 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09883 2297 1851 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09882 4478 1999 2297 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09881 544 549 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09880 4478 1591 549 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09879 549 581 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09878 229 222 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09877 4478 1591 222 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09876 222 238 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09875 2171 2656 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09874 1750 1590 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09873 4478 1782 1590 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09872 1590 1589 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09871 537 384 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09870 4478 1782 384 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09869 384 763 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09868 576 405 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09867 4478 1782 405 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09866 405 404 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09865 2655 2657 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09864 4478 2656 2657 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09863 2657 2695 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09862 2325 2357 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09861 2315 1415 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09860 4478 1421 2315 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09859 856 231 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09858 4478 1782 231 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09857 231 229 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09856 1107 2782 1108 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09855 4478 1126 1107 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09854 1111 1108 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09853 1882 2034 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_09852 2175 2924 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09851 2229 1893 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_09850 693 209 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09849 4478 207 209 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09848 209 1591 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09847 181 212 207 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09846 4478 210 181 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09845 521 1044 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09844 4478 828 747 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09843 747 826 746 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09842 746 825 827 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09841 1838 827 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09840 1109 1111 1115 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_09839 4478 1117 1109 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_09838 1975 1115 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09837 2783 2589 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09836 2600 2488 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09835 555 386 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09834 4478 385 386 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09833 386 401 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09832 1862 1503 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09831 4478 1589 1503 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09830 1503 1499 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09829 2513 2435 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_09828 1025 1564 1024 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09827 4478 1026 1025 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09826 1040 1024 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09825 2841 2481 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09824 4478 2423 2481 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09823 2481 2424 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09822 853 852 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09821 4478 2423 852 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09820 852 1704 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09819 765 764 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09818 4478 2423 764 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09817 764 1287 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09816 1669 1847 2002 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09815 4478 1709 1669 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09814 2694 2693 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09813 4478 2691 2693 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09812 2693 2695 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09811 332 294 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09810 4478 1782 294 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09809 294 291 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09808 2840 2698 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09807 4478 2696 2698 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09806 2698 2695 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09805 661 304 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09804 4478 1782 304 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09803 304 303 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09802 728 635 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09801 4478 1782 635 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09800 635 633 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09799 1472 1529 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09798 4478 1782 1529 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09797 1529 1527 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09796 2545 2781 2544 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09795 4478 2542 2545 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09794 291 241 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09793 4478 238 241 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09792 241 264 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09791 614 612 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09790 4478 605 612 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09789 612 608 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09788 1895 1780 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09787 4478 1785 1780 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09786 1780 1778 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09785 1785 1570 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09784 4478 1569 1570 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09783 1570 1572 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09782 1594 1591 1593 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09781 4478 1592 1594 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09780 1598 1593 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09779 2699 2323 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_09778 2123 2122 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09777 4478 2123 2124 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09776 2124 4350 2584 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09775 2271 2781 2457 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09774 4478 2390 2271 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09773 1599 1782 2447 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09772 4478 1598 1599 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09771 2360 1521 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09770 4478 1522 1521 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09769 1521 1458 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09768 784 785 2696 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09767 4478 783 784 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09766 2702 2120 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09765 4478 2118 2120 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09764 2120 2117 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09763 1455 1598 1911 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09762 4478 1460 1455 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09761 2227 805 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09760 4478 803 805 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09759 805 731 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09758 1470 1532 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09757 4478 1470 1469 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09756 1469 1468 2455 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09755 1457 1522 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09754 4478 1457 1459 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09753 1459 1458 2199 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09752 2114 2118 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09751 4478 2114 1969 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09750 1969 2117 2844 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09749 1041 1782 2435 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09748 4478 1040 1041 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09747 2429 2016 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09746 4478 2020 2016 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09745 2016 2022 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09744 1427 1782 1428 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09743 4478 1426 1427 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09742 1039 1040 2656 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09741 4478 1038 1039 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09740 2352 1596 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09739 4478 1754 1596 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09738 1596 1595 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09737 1320 1426 2357 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09736 4478 1319 1320 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09735 2021 2020 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09734 4478 2021 1956 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09733 1956 2022 2613 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09732 4478 367 364 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09731 366 1972 365 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09730 364 363 366 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09729 1423 1421 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09728 4478 1423 1422 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09727 1422 1420 1585 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09726 2808 2823 2809 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09725 4478 2930 2808 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09724 2815 2817 2814 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09723 4478 2937 2815 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09722 2824 2823 2825 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09721 4478 2937 2824 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09720 2933 2932 2934 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09719 4478 2937 2933 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09718 2323 2307 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09717 4478 2424 2323 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09716 742 823 829 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09715 4478 824 742 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09714 1850 2620 1999 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09713 4478 2111 1850 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09712 1417 2325 1421 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09711 4478 2111 1417 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09710 1597 2171 1754 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09709 4478 2111 1597 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09708 1955 2513 2020 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09707 4478 2111 1955 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09706 804 2222 803 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09705 4478 988 804 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09704 1968 2220 2118 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09703 4478 2111 1968 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09702 1461 2542 1522 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09701 4478 2111 1461 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09700 1467 2390 1532 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09699 4478 2111 1467 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09698 1564 367 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_09697 1835 1571 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09696 2423 1126 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09695 1591 520 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09694 1407 3226 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09693 2136 3905 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_09692 2284 3911 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09691 2778 3835 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09690 2937 2930 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_09689 785 703 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09688 4478 704 785 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09687 2390 2197 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_09686 1896 1526 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09685 4478 1527 1526 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09684 1526 1462 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09683 2217 1531 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09682 4478 1532 1531 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09681 1531 1465 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09680 1614 2070 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09679 1617 1621 1614 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09678 1615 1623 1617 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09677 1620 1623 1616 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09676 1616 1615 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09675 1619 1621 1620 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09674 1623 1622 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09673 4478 1623 1621 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09672 1618 1624 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09671 4478 1618 1619 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09670 4478 1617 2070 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09669 2070 1617 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09668 1615 1620 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09667 425 913 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09666 424 434 425 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09665 426 433 424 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09664 428 433 430 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09663 430 426 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09662 427 434 428 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09661 433 432 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09660 4478 433 434 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09659 429 435 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09658 4478 429 427 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09657 4478 424 913 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09656 913 424 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09655 426 428 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09654 193 723 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09653 310 317 193 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09652 309 321 310 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09651 312 321 192 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09650 192 309 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09649 194 317 312 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09648 321 314 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09647 4478 321 317 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09646 315 320 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09645 4478 315 194 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09644 4478 310 723 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09643 723 310 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09642 309 312 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09641 2207 2688 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09640 2208 2210 2207 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09639 2209 2216 2208 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09638 2213 2216 2206 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09637 2206 2209 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09636 2212 2210 2213 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09635 2216 2214 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09634 4478 2216 2210 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09633 2211 2215 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09632 4478 2211 2212 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09631 4478 2208 2688 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09630 2688 2208 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09629 2209 2213 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09628 4478 2192 2189 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09627 2192 2191 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09626 4478 2360 2193 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09625 2193 2195 2192 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09624 2182 2195 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09623 2183 2184 2182 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09622 2180 2190 2183 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09621 2187 2190 2181 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09620 2181 2180 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09619 2186 2184 2187 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09618 2190 2188 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09617 4478 2190 2184 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09616 2185 2189 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09615 4478 2185 2186 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09614 4478 2183 2195 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09613 2195 2183 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09612 2180 2187 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09611 4478 601 600 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09610 601 603 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09609 4478 2360 492 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09608 492 904 601 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09607 489 904 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09606 589 598 489 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09605 593 599 589 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09604 591 599 491 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09603 491 593 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09602 490 598 591 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09601 599 594 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09600 4478 599 598 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09599 597 600 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09598 4478 597 490 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09597 4478 589 904 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09596 904 589 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09595 593 591 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09594 4478 284 283 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09593 284 288 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09592 4478 2360 191 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09591 191 715 284 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09590 188 715 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09589 271 280 188 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09588 272 278 271 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09587 275 278 190 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09586 190 272 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09585 189 280 275 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09584 278 277 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09583 4478 278 280 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09582 274 283 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09581 4478 274 189 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09580 4478 271 715 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09579 715 271 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09578 272 275 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09577 4478 2363 2538 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09576 2363 2366 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09575 4478 2360 2267 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09574 2267 2826 2363 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09573 2536 2826 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09572 2535 2532 2536 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09571 2537 2533 2535 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09570 2534 2533 2540 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09569 2540 2537 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09568 2539 2532 2534 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09567 2533 2451 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09566 4478 2533 2532 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09565 2541 2538 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09564 4478 2541 2539 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09563 4478 2535 2826 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09562 2826 2535 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09561 2537 2534 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09560 4478 1643 1651 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09559 1643 1642 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09558 4478 2702 1644 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09557 1644 1812 1643 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09556 1649 1812 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09555 1650 1659 1649 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09554 1652 1658 1650 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09553 1654 1658 1655 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09552 1655 1652 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09551 1653 1659 1654 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09550 1658 1656 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09549 4478 1658 1659 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09548 1657 1651 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09547 4478 1657 1653 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09546 4478 1650 1812 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09545 1812 1650 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09544 1652 1654 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09543 1084 728 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09542 4478 763 1084 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09541 4478 1085 1082 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09540 1085 1084 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09539 4478 2702 1086 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09538 1086 1091 1085 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09537 1073 1091 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09536 1074 1080 1073 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09535 1075 1083 1074 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09534 1078 1083 1076 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09533 1076 1075 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09532 1079 1080 1078 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09531 1083 1081 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09530 4478 1083 1080 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09529 1077 1082 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09528 4478 1077 1079 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09527 4478 1074 1091 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09526 1091 1074 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09525 1075 1078 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09524 1379 661 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09523 4478 855 1379 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09522 4478 1380 1385 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09521 1380 1379 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09520 4478 2702 1381 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09519 1381 1382 1380 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09518 1383 1382 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09517 1384 1393 1383 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09516 1386 1394 1384 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09515 1389 1394 1388 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09514 1388 1386 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09513 1390 1393 1389 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09512 1394 1391 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09511 4478 1394 1393 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09510 1392 1385 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09509 4478 1392 1390 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09508 4478 1384 1382 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09507 1382 1384 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09506 1386 1389 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09505 2701 2699 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09504 4478 2840 2701 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09503 4478 2704 2708 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09502 2704 2701 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09501 4478 2702 2558 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09500 2558 2705 2704 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09499 2564 2705 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09498 2706 2715 2564 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09497 2709 2716 2706 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09496 2710 2716 2571 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09495 2571 2709 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09494 2570 2715 2710 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09493 2716 2713 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09492 4478 2716 2715 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09491 2714 2708 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09490 4478 2714 2570 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09489 4478 2706 2705 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09488 2705 2706 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09487 2709 2710 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09486 1641 1804 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09485 4478 1894 1641 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09484 4478 1639 1638 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09483 1639 1641 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09482 4478 2227 1640 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09481 1640 1810 1639 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09480 1629 1810 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09479 1630 1631 1629 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09478 1628 1637 1630 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09477 1635 1637 1634 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09476 1634 1628 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09475 1633 1631 1635 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09474 1637 1636 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09473 4478 1637 1631 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09472 1632 1638 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09471 4478 1632 1633 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09470 4478 1630 1810 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09469 1810 1630 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09468 1628 1635 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09467 452 658 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09466 4478 763 452 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09465 4478 453 455 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09464 453 452 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09463 4478 2227 454 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09462 454 1090 453 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09461 442 1090 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09460 444 451 442 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09459 445 449 444 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09458 447 449 446 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09457 446 445 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09456 443 451 447 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09455 449 448 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09454 4478 449 451 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09453 450 455 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09452 4478 450 443 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09451 4478 444 1090 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09450 1090 444 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09449 445 447 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09448 335 332 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09447 4478 855 335 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09446 4478 336 342 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09445 336 335 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09444 4478 2227 196 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09443 196 1371 336 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09442 197 1371 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09441 341 350 197 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09440 343 351 341 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09439 348 351 199 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09438 199 343 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09437 198 350 348 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09436 351 349 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09435 4478 351 350 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09434 352 342 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09433 4478 352 198 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09432 4478 341 1371 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09431 1371 341 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09430 343 348 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09429 2401 2699 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09428 4478 2694 2401 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09427 4478 2225 2233 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09426 2225 2401 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09425 4478 2227 2228 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09424 2228 2677 2225 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09423 2231 2677 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09422 2232 2241 2231 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09421 2234 2240 2232 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09420 2237 2240 2236 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09419 2236 2234 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09418 2235 2241 2237 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09417 2240 2238 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09416 4478 2240 2241 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09415 2239 2233 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09414 4478 2239 2235 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09413 4478 2232 2677 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09412 2677 2232 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09411 2234 2237 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09410 2096 1896 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09409 4478 2002 2096 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09408 4478 2097 2106 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09407 2097 2096 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09406 4478 2099 1964 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09405 1964 2455 2097 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09404 1965 2099 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09403 2104 2108 1965 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09402 2101 2112 2104 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09401 2103 2112 1966 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09400 1966 2101 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09399 1967 2108 2103 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09398 2112 2105 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09397 4478 2112 2108 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09396 2107 2106 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09395 4478 2107 1967 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09394 4478 2104 2099 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09393 2099 2104 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09392 2101 2103 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09391 649 441 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09390 4478 765 649 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09389 4478 653 651 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09388 653 649 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09387 4478 926 500 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09386 500 2455 653 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09385 497 926 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09384 637 646 497 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09383 640 647 637 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09382 641 647 499 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09381 499 640 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09380 498 646 641 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09379 647 644 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09378 4478 647 646 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09377 648 651 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09376 4478 648 498 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09375 4478 637 926 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09374 926 637 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09373 640 641 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09372 654 328 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09371 4478 853 654 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09370 4478 657 796 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09369 657 654 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09368 4478 1206 501 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09367 501 2455 657 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09366 790 1206 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09365 791 787 790 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09364 794 788 791 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09363 792 788 795 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09362 795 794 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09361 793 787 792 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09360 788 726 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09359 4478 788 787 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09358 799 796 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09357 4478 799 793 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09356 4478 791 1206 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09355 1206 791 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09354 794 792 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09353 2459 2457 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09352 4478 2841 2459 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09351 4478 2555 2556 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09350 2555 2459 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09349 4478 2684 2456 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09348 2456 2455 2555 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09347 2547 2684 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09346 2552 2546 2547 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09345 2551 2548 2552 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09344 2549 2548 2550 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09343 2550 2551 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09342 2553 2546 2549 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09341 2548 2454 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09340 4478 2548 2546 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09339 2554 2556 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09338 4478 2554 2553 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09337 4478 2552 2684 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09336 2684 2552 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09335 2551 2549 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09334 1897 1895 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09333 4478 2002 1897 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09332 4478 1899 1906 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09331 1899 1897 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09330 4478 2065 1898 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09329 1898 2199 1899 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09328 1900 2065 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09327 1902 1910 1900 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09326 1903 1909 1902 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09325 1905 1909 1904 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09324 1904 1903 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09323 1901 1910 1905 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09322 1909 1907 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09321 4478 1909 1910 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09320 1908 1906 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09319 4478 1908 1901 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09318 4478 1902 2065 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09317 2065 1902 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09316 1903 1905 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09315 630 614 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09314 4478 765 630 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09313 4478 632 626 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09312 632 630 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09311 4478 1063 496 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09310 496 2199 632 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09309 493 1063 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09308 617 624 493 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09307 616 627 617 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09306 622 627 495 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09305 495 616 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09304 494 624 622 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09303 627 625 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09302 4478 627 624 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09301 620 626 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09300 4478 620 494 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09299 4478 617 1063 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09298 1063 617 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09297 616 622 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09296 1200 296 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09295 4478 853 1200 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09294 4478 1201 1363 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09293 1201 1200 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09292 4478 1357 1071 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09291 1071 2199 1201 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09290 1356 1357 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09289 1361 1366 1356 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09288 1358 1367 1361 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09287 1360 1367 1359 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09286 1359 1358 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09285 1365 1366 1360 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09284 1367 1362 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09283 4478 1367 1366 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09282 1364 1363 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09281 4478 1364 1365 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09280 4478 1361 1357 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09279 1357 1361 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09278 1358 1360 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09277 2453 2544 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09276 4478 2841 2453 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09275 4478 2200 2372 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09274 2200 2453 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09273 4478 2664 2201 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09272 2201 2199 2200 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09271 2268 2664 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09270 2370 2379 2268 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09269 2373 2380 2370 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09268 2377 2380 2270 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09267 2270 2373 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09266 2269 2379 2377 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09265 2380 2378 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09264 4478 2380 2379 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09263 2374 2372 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09262 4478 2374 2269 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09261 4478 2370 2664 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09260 2664 2370 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09259 2373 2377 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09258 1474 1472 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09257 4478 2002 1474 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09256 4478 1539 1478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09255 1539 1474 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09254 4478 1915 1475 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09253 1475 2844 1539 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09252 1387 1915 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09251 1541 1485 1387 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09250 1543 1486 1541 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09249 1542 1486 1480 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09248 1480 1543 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09247 1479 1485 1542 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09246 1486 1484 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09245 4478 1486 1485 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09244 1483 1478 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09243 4478 1483 1479 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09242 4478 1541 1915 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09241 1915 1541 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09240 1543 1542 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09239 934 728 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09238 4478 765 934 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09237 4478 935 943 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09236 935 934 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09235 4478 1092 802 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09234 802 2844 935 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09233 811 1092 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09232 941 950 811 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09231 944 951 941 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09230 945 951 817 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09229 817 944 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09228 816 950 945 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09227 951 948 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09226 4478 951 950 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09225 949 943 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09224 4478 949 816 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09223 4478 941 1092 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09222 1092 941 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09221 944 945 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09220 937 661 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09219 4478 853 937 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09218 4478 940 938 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09217 940 937 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09216 4478 1226 806 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09215 806 2844 940 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09214 810 1226 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09213 809 807 810 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09212 812 808 809 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09211 813 808 814 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09210 814 812 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09209 815 807 813 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09208 808 733 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09207 4478 808 807 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09206 818 938 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09205 4478 818 815 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09204 4478 809 1226 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09203 1226 809 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09202 812 813 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09201 2842 2840 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09200 4478 2841 2842 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09199 4478 2843 2850 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09198 2843 2842 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09197 4478 2846 2845 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09196 2845 2844 2843 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09195 2847 2846 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09194 2848 2856 2847 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09193 2849 2857 2848 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09192 2853 2857 2852 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09191 2852 2849 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09190 2851 2856 2853 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09189 2857 2854 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09188 4478 2857 2856 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09187 2855 2850 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09186 4478 2855 2851 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09185 4478 2848 2846 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09184 2846 2848 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09183 2849 2853 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09182 1925 1804 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09181 4478 2002 1925 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09180 4478 1926 1931 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09179 1926 1925 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09178 4478 1928 1927 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09177 1927 2463 1926 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09176 1929 1928 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09175 1930 1938 1929 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09174 1932 1937 1930 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09173 1935 1937 1934 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09172 1934 1932 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09171 1933 1938 1935 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09170 1937 1936 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09169 4478 1937 1938 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09168 1939 1931 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09167 4478 1939 1933 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09166 4478 1930 1928 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09165 1928 1930 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09164 1932 1935 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09163 662 658 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09162 4478 765 662 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09161 4478 665 669 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09160 665 662 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09159 4478 1095 502 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09158 502 730 665 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09157 503 1095 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09156 667 677 503 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09155 670 678 667 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09154 673 678 505 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09153 505 670 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09152 504 677 673 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09151 678 676 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09150 4478 678 677 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09149 679 669 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09148 4478 679 504 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09147 4478 667 1095 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09146 1095 667 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09145 670 673 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09144 458 332 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09143 4478 853 458 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09142 4478 461 464 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09141 461 458 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09140 4478 1232 460 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09139 460 730 461 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09138 462 1232 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09137 463 472 462 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09136 465 471 463 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09135 468 471 467 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09134 467 465 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09133 466 472 468 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09132 471 469 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09131 4478 471 472 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09130 470 464 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09129 4478 470 466 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09128 4478 463 1232 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09127 1232 463 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09126 465 468 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09125 2462 2694 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09124 4478 2841 2462 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09123 4478 2557 2566 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09122 2557 2462 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09121 4478 2561 2464 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09120 2464 2463 2557 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09119 2563 2561 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09118 2562 2559 2563 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09117 2565 2560 2562 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09116 2567 2560 2568 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09115 2568 2565 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09114 2569 2559 2567 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09113 2560 2465 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09112 4478 2560 2559 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09111 2572 2566 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09110 4478 2572 2569 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09109 4478 2562 2561 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09108 2561 2562 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09107 2565 2567 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09106 4478 1512 1440 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09105 1512 1438 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09104 4478 1441 1439 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09103 1439 2635 1512 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09102 1438 576 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09101 4478 853 1438 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09100 1019 1298 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09099 1128 1136 1019 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09098 1129 1137 1128 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09097 1130 1137 1022 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09096 1022 1129 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09095 1023 1136 1130 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09094 1137 1134 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09093 4478 1137 1136 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09092 1135 1133 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09091 4478 1135 1023 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09090 4478 1128 1298 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09089 1298 1128 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09088 1129 1130 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09087 1867 2023 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09086 1869 1877 1867 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09085 1868 1876 1869 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09084 1874 1876 1873 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09083 1873 1868 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09082 1871 1877 1874 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09081 1876 1875 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09080 4478 1876 1877 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09079 1872 1870 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09078 4478 1872 1871 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09077 4478 1869 2023 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09076 2023 1869 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09075 1868 1874 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09074 4478 1752 1870 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09073 1752 1751 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09072 4478 2023 1678 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09071 1678 2635 1752 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09070 1751 1750 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09069 4478 2002 1751 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09068 2755 2806 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09067 2756 2765 2755 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09066 2757 2762 2756 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09065 2759 2762 2758 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09064 2758 2757 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09063 2764 2765 2759 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09062 2762 2760 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09061 4478 2762 2765 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09060 2763 2761 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09059 4478 2763 2764 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09058 4478 2756 2806 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09057 2806 2756 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09056 2757 2759 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09055 4478 2479 2482 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09054 2483 2806 2482 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09053 2482 3911 2483 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09052 2489 2488 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09051 2490 2485 2489 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09050 2491 2486 2490 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09049 2487 2486 2493 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09048 2493 2491 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09047 2492 2485 2487 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09046 2486 2427 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09045 4478 2486 2485 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09044 2494 2594 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09043 4478 2494 2492 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09042 4478 2490 2488 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09041 2488 2490 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09040 2491 2487 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09039 4478 2141 2147 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09038 2141 2140 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09037 4478 2139 2142 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09036 2142 3911 2141 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_09035 2140 2138 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_09034 1010 1032 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09033 1012 1014 1010 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09032 1011 1021 1012 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09031 1016 1021 1018 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09030 1018 1011 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09029 1017 1014 1016 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09028 1021 1020 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09027 4478 1021 1014 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09026 1015 1013 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09025 4478 1015 1017 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09024 4478 1012 1032 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09023 1032 1012 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09022 1011 1016 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09021 1001 1412 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_09020 1947 2055 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09019 1988 1996 1947 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09018 1990 1997 1988 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09017 1993 1997 1949 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09016 1949 1990 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09015 1948 1996 1993 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09014 1997 1995 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09013 4478 1997 1996 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09012 1998 2005 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09011 4478 1998 1948 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09010 4478 1988 2055 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09009 2055 1988 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09008 1990 1993 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09007 2005 2008 1951 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09006 1950 2003 2005 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_09005 4478 2002 1951 4478 tp L=0.32U W=4.05U AS=3.0375P AD=3.0375P PS=9.6U PD=9.6U 
Mtr_09004 1951 2004 4478 4478 tp L=0.32U W=4.05U AS=3.0375P AD=3.0375P PS=9.6U PD=9.6U 
Mtr_09003 1951 2001 1950 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_09002 2003 1999 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_09001 2504 2801 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_09000 2604 2610 2504 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08999 2605 2611 2604 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08998 2607 2611 2508 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08997 2508 2605 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08996 2509 2610 2607 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08995 2611 2609 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08994 4478 2611 2610 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08993 2612 2614 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08992 4478 2612 2509 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08991 4478 2604 2801 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08990 2801 2604 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08989 2605 2607 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08988 4478 2615 2614 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08987 2615 2619 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08986 4478 2801 2512 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08985 2512 2613 2615 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08984 2619 2617 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08983 4478 2841 2619 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08982 485 1326 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08981 564 569 485 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08980 563 567 564 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08979 561 567 487 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08978 487 563 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08977 486 569 561 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08976 567 566 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08975 4478 567 569 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08974 568 573 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08973 4478 568 486 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08972 4478 564 1326 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08971 1326 564 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08970 563 561 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08969 2012 1862 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08968 4478 1894 2012 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08967 4478 2015 2153 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08966 2015 2012 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08965 4478 2429 1954 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08964 1954 2161 2015 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08963 2152 2161 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08962 2151 2154 2152 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08961 2149 2159 2151 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08960 2157 2159 2150 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08959 2150 2149 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08958 2156 2154 2157 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08957 2159 2158 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08956 4478 2159 2154 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08955 2155 2153 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08954 4478 2155 2156 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08953 4478 2151 2161 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08952 2161 2151 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08951 2149 2157 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08950 553 555 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08949 4478 763 553 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08948 4478 550 547 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08947 550 553 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08946 4478 2429 484 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08945 484 1160 550 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08944 480 1160 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08943 529 535 480 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08942 528 536 529 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08941 527 536 482 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08940 482 528 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08939 481 535 527 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08938 536 531 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08937 4478 536 535 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08936 533 547 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08935 4478 533 481 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08934 4478 529 1160 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08933 1160 529 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08932 528 527 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08931 400 402 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08930 4478 855 400 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08929 4478 398 397 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08928 398 400 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08927 4478 2429 399 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08926 399 1152 398 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08925 387 1152 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08924 388 395 387 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08923 389 396 388 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08922 391 396 390 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08921 390 389 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08920 394 395 391 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08919 396 392 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08918 4478 396 395 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08917 393 397 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08916 4478 393 394 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08915 4478 388 1152 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08914 1152 388 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08913 389 391 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08912 2432 2699 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08911 4478 2617 2432 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08910 4478 2510 2511 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08909 2510 2432 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08908 4478 2429 2430 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08907 2430 2497 2510 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08906 2501 2497 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08905 2502 2498 2501 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08904 2503 2499 2502 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08903 2500 2499 2506 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08902 2506 2503 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08901 2505 2498 2500 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08900 2499 2428 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08899 4478 2499 2498 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08898 2507 2511 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08897 4478 2507 2505 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08896 4478 2502 2497 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08895 2497 2502 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08894 2503 2500 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08893 1567 1708 1718 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08892 1718 2297 1567 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08891 4478 2004 1567 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08890 1567 1894 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08889 1670 1878 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08888 1716 1727 1670 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08887 1719 1728 1716 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08886 1723 1728 1672 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08885 1672 1719 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08884 1671 1727 1723 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08883 1728 1726 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08882 4478 1728 1727 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08881 1722 1718 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08880 4478 1722 1671 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08879 4478 1716 1878 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08878 1878 1716 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08877 1719 1723 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08876 754 877 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08875 836 842 754 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08874 835 844 836 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08873 837 844 759 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08872 759 835 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08871 760 842 837 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08870 844 839 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08869 4478 844 842 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08868 840 845 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08867 4478 840 760 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08866 4478 836 877 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08865 877 836 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08864 835 837 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08863 368 708 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08862 369 377 368 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08861 370 378 369 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08860 374 378 373 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08859 373 370 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08858 371 377 374 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08857 378 376 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08856 4478 378 377 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08855 372 380 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08854 4478 372 371 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08853 4478 369 708 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08852 708 369 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08851 370 374 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08850 2767 2802 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08849 2771 2776 2767 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08848 2772 2777 2771 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08847 2768 2777 2770 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08846 2770 2772 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08845 2769 2776 2768 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08844 2777 2773 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08843 4478 2777 2776 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08842 2775 2774 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08841 4478 2775 2769 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08840 4478 2771 2802 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08839 2802 2771 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08838 2772 2768 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08837 1600 1750 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08836 4478 1894 1600 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08835 4478 1601 1608 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08834 1601 1600 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08833 4478 2352 1602 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08832 1602 1886 1601 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08831 1603 1886 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08830 1607 1612 1603 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08829 1604 1613 1607 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08828 1606 1613 1605 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08827 1605 1604 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08826 1611 1612 1606 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08825 1613 1609 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08824 4478 1613 1612 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08823 1610 1608 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08822 4478 1610 1611 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08821 4478 1607 1886 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08820 1886 1607 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08819 1604 1606 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08818 255 385 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08817 4478 537 255 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08816 4478 257 258 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08815 257 255 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08814 4478 1170 187 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08813 187 1061 257 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08812 184 1061 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08811 248 253 184 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08810 247 250 248 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08809 245 250 186 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08808 186 247 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08807 185 253 245 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08806 250 249 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08805 4478 250 253 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08804 251 258 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08803 4478 251 185 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08802 4478 248 1061 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08801 1061 248 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08800 247 245 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08799 409 576 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08798 4478 855 409 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08797 4478 410 416 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08796 410 409 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08795 4478 1170 411 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08794 411 1348 410 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08793 414 1348 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08792 415 417 414 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08791 412 422 415 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08790 420 422 413 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08789 413 412 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08788 419 417 420 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08787 422 421 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08786 4478 422 417 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08785 418 416 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08784 4478 418 419 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08783 4478 415 1348 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08782 1348 415 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08781 412 420 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08780 2641 2699 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08779 4478 2655 2641 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08778 4478 2353 2647 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08777 2353 2641 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08776 4478 2352 2266 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08775 2266 2643 2353 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08774 2528 2643 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08773 2646 2648 2528 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08772 2645 2654 2646 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08771 2651 2654 2530 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08770 2530 2645 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08769 2531 2648 2651 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08768 2654 2653 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08767 4478 2654 2648 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08766 2649 2647 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08765 4478 2649 2531 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08764 4478 2646 2643 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08763 2643 2646 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08762 2645 2651 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08761 1673 1747 1738 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08760 1738 2315 1673 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08759 4478 1730 1673 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08758 1673 1894 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08757 1674 1885 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08756 1737 1743 1674 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08755 1736 1745 1737 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08754 1741 1745 1676 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08753 1676 1736 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08752 1675 1743 1741 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08751 1745 1744 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08750 4478 1745 1743 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08749 1739 1738 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08748 4478 1739 1675 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08747 4478 1737 1885 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08746 1885 1737 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08745 1736 1741 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08744 483 696 755 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08743 755 2315 483 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08742 4478 544 483 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08741 483 537 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08740 752 1051 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08739 753 748 752 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08738 751 749 753 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08737 750 749 757 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08736 757 751 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08735 756 748 750 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08734 749 695 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08733 4478 749 748 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08732 758 755 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08731 4478 758 756 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08730 4478 753 1051 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08729 1051 753 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08728 751 750 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08727 775 859 867 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08726 867 2315 775 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08725 4478 856 775 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08724 775 855 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08723 778 1347 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08722 861 869 778 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08721 862 870 861 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08720 864 870 779 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08719 779 862 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08718 780 869 864 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08717 870 866 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08716 4478 870 869 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08715 868 867 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08714 4478 868 780 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08713 4478 861 1347 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08712 1347 861 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08711 862 864 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08710 2253 2356 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08709 2305 2309 2253 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08708 2303 2313 2305 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08707 2311 2313 2252 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08706 2252 2303 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08705 2254 2309 2311 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08704 2313 2312 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08703 4478 2313 2309 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08702 2308 2317 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08701 4478 2308 2254 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08700 4478 2305 2356 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08699 2356 2305 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08698 2303 2311 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08697 1863 1862 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08696 4478 2002 1863 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08695 4478 1866 1865 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08694 1866 1863 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08693 4478 2027 1864 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08692 1864 2613 1866 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08691 1853 2027 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08690 1852 1860 1853 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08689 1854 1861 1852 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08688 1857 1861 1858 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08687 1858 1854 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08686 1855 1860 1857 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08685 1861 1859 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08684 4478 1861 1860 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08683 1856 1865 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08682 4478 1856 1855 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08681 4478 1852 2027 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08680 2027 1852 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08679 1854 1857 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08678 701 555 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08677 4478 765 701 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08676 4478 776 777 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08675 776 701 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08674 4478 1030 702 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08673 702 2613 776 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08672 770 1030 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08671 771 766 770 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08670 769 767 771 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08669 768 767 773 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08668 773 769 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08667 772 766 768 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08666 767 700 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08665 4478 767 766 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08664 774 777 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08663 4478 774 772 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08662 4478 771 1030 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08661 1030 771 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08660 769 768 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08659 572 402 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08658 4478 853 572 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08657 4478 574 573 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08656 574 572 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08655 4478 1326 488 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08654 488 2613 574 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08653 4478 2497 2445 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08652 2445 2435 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08651 2445 2438 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08650 4478 2450 2524 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08649 2526 2524 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08648 4478 2439 2524 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08647 2524 2440 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08646 4478 2643 2439 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08645 2439 2656 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08644 2439 2438 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08643 4478 2802 2440 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08642 2440 2437 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08641 2440 2438 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08640 4478 2688 2450 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08639 2450 2197 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08638 2450 2198 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08637 1354 1352 1355 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_08636 4478 1353 1354 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_08635 3111 1355 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08634 4478 1351 1353 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08633 1353 1372 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08632 4478 1350 1353 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08631 1353 1368 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08630 4478 1382 1368 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08629 1368 2696 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08628 1368 1376 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08627 4478 1347 1351 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08626 1351 2357 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08625 1351 1349 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08624 4478 1371 1372 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08623 1372 1911 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08622 1372 1376 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08621 4478 1348 1350 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08620 1350 2656 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08619 1350 1349 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08618 4478 1180 1352 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08617 1352 1214 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08616 4478 1179 1352 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08615 1352 1331 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08614 1333 2488 1331 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08613 1333 1328 1332 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08612 1332 1329 1333 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08611 1332 1326 1327 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08610 4478 1337 1327 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08609 1331 1330 1333 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08608 1327 1441 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08607 1327 1445 1332 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08606 1335 2171 1337 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08605 4478 1334 1335 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08604 1443 2513 1445 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08603 4478 1442 1443 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08602 1322 2325 1329 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08601 4478 1323 1322 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08600 1325 2620 1330 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08599 4478 1323 1325 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08598 1143 1152 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_08597 1212 1232 1214 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08596 1212 1206 1209 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08595 1209 1207 1212 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08594 1209 1226 1208 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08593 4478 1357 1208 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08592 1214 1219 1212 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08591 1208 1369 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08590 1208 1216 1209 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08589 1370 2542 1369 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08588 4478 1376 1370 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08587 1215 2220 1216 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08586 4478 1217 1215 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08585 1203 2390 1207 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08584 4478 1204 1203 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08583 1218 2222 1219 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08582 4478 1217 1218 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08581 4478 709 781 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08580 1179 781 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08579 4478 713 781 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08578 781 710 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08577 4478 723 713 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08576 713 2197 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08575 713 714 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08574 4478 708 710 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08573 710 1428 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08572 710 714 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08571 4478 715 709 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08570 709 2447 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08569 709 714 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08568 1059 1057 1060 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_08567 4478 1058 1059 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_08566 3377 1060 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08565 4478 1055 1058 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08564 1058 1056 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08563 4478 1066 1058 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08562 1058 1070 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08561 4478 1091 1070 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08560 1070 2696 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08559 1070 1072 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08558 1055 1166 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08557 4478 1298 1055 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08556 1165 2171 1166 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08555 4478 1164 1165 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08554 4478 1051 1056 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08553 1056 2357 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08552 1056 1052 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08551 4478 1037 1057 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08550 1057 898 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08549 4478 892 1057 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08548 1057 930 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08547 800 1095 930 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08546 800 926 797 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08545 797 1088 800 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08544 797 1092 798 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08543 4478 1063 798 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08542 930 929 800 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08541 798 1377 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08540 798 933 797 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08539 1378 2542 1377 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08538 4478 1376 1378 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08537 801 2220 933 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08536 4478 932 801 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08535 1089 2390 1088 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08534 4478 1087 1089 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08533 789 2222 929 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08532 4478 924 789 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08531 1036 1032 1037 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08530 1037 1035 1036 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08529 1036 1033 1034 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08528 1034 1044 1036 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08527 4478 1030 1034 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08526 1034 1147 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08525 1146 2513 1147 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08524 4478 1145 1146 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08523 1029 2325 1033 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08522 4478 1027 1029 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08521 1031 2620 1035 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08520 4478 1027 1031 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08519 4478 888 890 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08518 892 890 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08517 4478 1062 890 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08516 890 887 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08515 2205 2203 2204 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_08514 4478 2202 2205 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_08513 3118 2204 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08512 1959 2168 2044 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08511 1959 2027 1960 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08510 1960 2031 1959 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08509 1960 2023 1958 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08508 4478 2055 1958 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08507 2044 2026 1959 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08506 1958 2165 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08505 1958 2033 1960 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08504 2163 2620 2165 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08503 4478 2166 2163 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08502 1962 2171 2033 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08501 4478 2032 1962 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08500 2160 2161 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_08499 1918 1928 2042 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08498 1918 2099 1917 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08497 1917 1914 1918 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08496 1917 1915 1916 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08495 4478 2065 1916 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08494 2042 1923 1918 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08493 1916 1920 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08492 1916 2094 1917 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08491 4478 2179 2040 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08490 2043 2040 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08489 4478 2064 2040 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08488 2040 2035 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08487 2127 2516 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08486 2128 2134 2127 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08485 2129 2135 2128 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08484 2126 2135 2125 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08483 2125 2129 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08482 2133 2134 2126 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08481 2135 2131 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08480 4478 2135 2134 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08479 2132 2130 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08478 4478 2132 2133 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08477 4478 2128 2516 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08476 2516 2128 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08475 2129 2126 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08474 1305 1328 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08473 1306 1313 1305 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08472 1307 1316 1306 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08471 1308 1316 1309 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08470 1309 1307 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08469 1314 1313 1308 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08468 1316 1310 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08467 4478 1316 1313 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08466 1312 1311 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08465 4478 1312 1314 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08464 4478 1306 1328 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08463 1328 1306 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08462 1307 1308 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08461 4478 1139 1311 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08460 1139 1138 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08459 4478 1328 1028 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08458 1028 1585 1139 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08457 1138 856 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08456 4478 853 1138 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08455 354 1044 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08454 353 362 354 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08453 356 360 353 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08452 358 360 357 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08451 357 356 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08450 355 362 358 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08449 360 359 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08448 4478 360 362 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08447 361 511 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08446 4478 361 355 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08445 4478 353 1044 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08444 1044 353 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08443 356 358 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08442 511 513 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08441 477 1044 476 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08440 477 743 4478 4478 tp L=0.35U W=4.05U AS=3.1185P AD=3.1185P PS=9.65U PD=9.65U 
Mtr_08439 4478 516 477 4478 tp L=0.35U W=4.05U AS=3.1185P AD=3.1185P PS=9.65U PD=9.65U 
Mtr_08438 476 510 513 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08437 513 745 477 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08436 1574 2168 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08435 1576 1583 1574 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08434 1575 1584 1576 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08433 1579 1584 1578 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08432 1578 1575 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08431 1580 1583 1579 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08430 1584 1581 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08429 4478 1584 1583 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08428 1577 1582 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08427 4478 1577 1580 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08426 4478 1576 2168 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08425 2168 1576 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08424 1575 1579 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08423 4478 1586 1582 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08422 1586 1588 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08421 4478 2168 1587 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08420 1587 1585 1586 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08419 1588 1730 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08418 4478 2002 1588 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08417 2521 2636 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08416 2626 2633 2521 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08415 2625 2630 2626 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08414 2628 2630 2522 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08413 2522 2625 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08412 2523 2633 2628 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08411 2630 2629 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08410 4478 2630 2633 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08409 2631 2634 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08408 4478 2631 2523 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08407 4478 2626 2636 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08406 2636 2626 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08405 2625 2628 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08404 4478 2638 2634 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08403 2638 2639 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08402 4478 2636 2525 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08401 2525 2635 2638 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08400 2639 2655 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08399 4478 2841 2639 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08398 1324 1441 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08397 1507 1436 1324 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08396 1509 1437 1507 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08395 1510 1437 1431 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08394 1431 1509 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08393 1430 1436 1510 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08392 1437 1434 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08391 4478 1437 1436 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08390 1435 1440 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08389 4478 1435 1430 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08388 4478 1507 1441 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08387 1441 1507 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08386 1509 1510 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08385 4478 1156 1158 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08384 1184 1328 1158 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08383 1158 1339 1184 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08382 1340 2335 1339 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08381 4478 1341 1340 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08380 4478 2924 1154 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08379 1156 1154 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08378 4478 1159 1154 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08377 1154 1152 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08376 4478 1067 3380 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08375 3380 1068 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08374 3380 1069 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08373 1069 911 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08372 911 907 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08371 4478 914 911 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08370 911 908 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08369 4478 921 911 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08368 4478 904 907 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08367 907 1893 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08366 907 920 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08365 4478 913 914 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08364 914 2934 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08363 914 920 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08362 4478 1032 908 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08361 908 2812 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08360 908 884 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08359 4478 926 921 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08358 921 2825 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08357 921 920 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08356 1097 1095 1096 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08355 1097 1091 1094 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08354 1094 1221 1097 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08353 1094 1092 1093 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08352 4478 1090 1093 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08351 1096 1374 1097 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08350 1093 1098 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08349 1093 1103 1094 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08348 1099 2229 1098 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08347 4478 1101 1099 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08346 1102 2414 1103 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08345 4478 1101 1102 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08344 1220 1646 1221 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08343 4478 1222 1220 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08342 1375 2410 1374 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08341 4478 1373 1375 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08340 4478 877 871 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08339 871 706 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08338 871 707 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08337 4478 1030 874 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08336 874 2809 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08335 874 884 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08334 4478 1169 1054 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08333 1068 1054 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08332 4478 1064 1054 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08331 1054 1053 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08330 4478 1063 1064 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08329 1064 2814 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08328 1064 1065 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08327 1047 1044 1053 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08326 1053 1049 1047 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08325 1047 1045 1046 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08324 1046 1051 1047 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08323 4478 1061 1046 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08322 1046 1338 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08321 1336 2175 1338 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08320 4478 1341 1336 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08319 1043 1882 1045 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08318 4478 1042 1043 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08317 1050 2335 1049 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08316 4478 1048 1050 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08315 4478 1167 1171 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08314 1169 1298 1171 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08313 1171 1449 1169 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08312 1448 2337 1449 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08311 4478 1452 1448 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08310 4478 2924 1163 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08309 1167 1163 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08308 4478 1159 1163 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08307 1163 1160 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08306 4478 2087 3221 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08305 3221 2088 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08304 3221 2092 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08303 4478 2195 2196 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08302 2196 2827 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08301 2196 2194 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08300 4478 2070 2076 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08299 2076 2934 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08298 2076 2081 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08297 4478 2055 2075 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08296 2075 2812 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08295 2075 2081 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08294 4478 2099 2084 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08293 2084 2825 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08292 2084 2081 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08291 1685 1928 1815 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08290 1685 1812 1684 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08289 1684 1813 1685 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08288 1684 1915 1683 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08287 4478 1810 1683 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08286 1815 1821 1685 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08285 1683 1819 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08284 1683 1825 1684 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08283 1686 2229 1819 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08282 4478 1824 1686 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08281 1688 2414 1825 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08280 4478 1824 1688 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08279 1645 1646 1813 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08278 4478 1647 1645 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08277 1687 2410 1821 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08276 4478 1824 1687 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08275 4478 1878 1764 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08274 1764 2034 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08273 1764 1770 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08272 4478 2027 1765 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08271 1765 2809 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08270 1765 1770 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08269 4478 2170 2054 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08268 2088 2054 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08267 4478 2066 2054 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08266 2054 2050 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08265 4478 2065 2066 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08264 2066 2814 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08263 2066 2081 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08262 1889 2023 2050 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08261 2050 1891 1889 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08260 1889 1887 1888 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08259 1888 1886 1889 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08258 4478 1885 1888 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08257 1888 1884 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08256 1880 1882 1884 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08255 4478 1881 1880 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08254 1680 2175 1887 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08253 4478 1770 1680 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08252 1890 2337 1891 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08251 4478 1892 1890 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08250 4478 2167 2169 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08249 2170 2168 2169 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08248 2169 2173 2170 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08247 2174 2335 2173 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08246 4478 2172 2174 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08245 4478 2924 2162 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08244 2167 2162 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08243 4478 2172 2162 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08242 2162 2161 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08241 2543 2668 2669 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_08240 4478 2676 2543 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_08239 3289 2669 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08238 4478 2672 2676 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08237 2676 2670 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08236 4478 2680 2676 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08235 2676 2671 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08234 4478 2705 2671 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08233 2671 2696 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08232 2671 2460 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08231 2672 2622 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08230 4478 2806 2672 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08229 2515 2620 2622 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08228 4478 2621 2515 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08227 4478 2356 2670 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08226 2670 2357 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08225 2670 2355 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08224 4478 2677 2680 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08223 2680 2691 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08222 2680 2683 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08221 4478 2444 2668 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08220 2668 2529 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08219 4478 2526 2668 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08218 2668 2443 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08217 2274 2561 2443 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08216 2274 2684 2273 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08215 2273 2392 2274 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08214 2273 2846 2272 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08213 4478 2664 2272 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08212 2443 2388 2274 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08211 2272 2394 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08210 2272 2384 2273 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08209 2276 2542 2394 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08208 4478 2395 2276 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08207 2221 2220 2384 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08206 4478 2223 2221 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08205 2275 2390 2392 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08204 4478 2391 2275 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08203 2224 2222 2388 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08202 4478 2223 2224 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08201 2260 2516 2444 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08200 2444 2327 2260 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08199 2260 2328 2259 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08198 2259 2636 2260 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08197 4478 2801 2259 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08196 2259 2332 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08195 2261 2513 2332 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08194 4478 2334 2261 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08193 2164 2171 2328 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08192 4478 2166 2164 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08191 2258 2325 2327 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08190 4478 2324 2258 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08189 4478 2826 2449 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08188 2449 2447 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08187 2449 2448 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08186 4478 1558 1560 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08185 1560 1558 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08184 4478 1558 1560 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08183 1558 1559 1557 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08182 4478 1563 1558 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08181 1559 1563 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08180 1560 1558 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08179 1558 3226 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08178 1562 1972 1563 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08177 4478 1561 1562 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08176 4478 3229 3230 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08175 3230 3229 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08174 4478 3229 3230 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08173 3229 3228 3297 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08172 4478 3232 3229 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08171 3228 3232 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08170 3230 3229 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08169 3229 3835 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08168 3232 3298 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08167 4478 3299 3298 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08166 3298 3233 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08165 4478 2839 3560 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08164 3560 2834 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08163 3560 2835 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08162 2835 2833 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08161 2833 2832 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08160 4478 2829 2833 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08159 2833 2830 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08158 4478 2831 2833 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08157 4478 2826 2832 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08156 2832 2827 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08155 2832 2828 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08154 4478 2688 2829 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08153 2829 2934 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08152 2829 2687 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08151 4478 2806 2830 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08150 2830 2812 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08149 2830 2807 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08148 4478 2684 2831 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08147 2831 2825 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08146 2831 2687 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08145 2839 2838 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08144 4478 2836 2838 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08143 2838 2837 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08142 2279 2561 2837 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08141 2279 2705 2278 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08140 2278 2404 2279 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08139 2278 2846 2277 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08138 4478 2677 2277 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08137 2837 2411 2279 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08136 2277 2402 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08135 2277 2416 2278 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08134 2230 2229 2402 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08133 4478 2226 2230 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08132 2281 2414 2416 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08131 4478 2415 2281 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08130 1648 1646 2404 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08129 4478 1647 1648 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08128 2280 2410 2411 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08127 4478 2415 2280 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08126 2836 2805 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08125 4478 2803 2805 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08124 2805 2804 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08123 4478 2802 2804 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08122 2804 2811 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08121 2804 2807 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08120 4478 2801 2803 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08119 2803 2809 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08118 2803 2807 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08117 4478 2660 2661 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08116 2834 2661 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08115 4478 2665 2661 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08114 2661 2659 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08113 4478 2664 2665 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08112 2665 2814 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08111 2665 2682 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08110 2264 2636 2659 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08109 2659 2346 2264 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08108 2264 2345 2265 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08107 2265 2643 2264 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08106 4478 2356 2265 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08105 2265 2341 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08104 1883 1882 2341 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08103 4478 1881 1883 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08102 2177 2175 2345 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08101 4478 2176 2177 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08100 2263 2337 2346 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08099 4478 2338 2263 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08098 4478 2520 2518 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08097 2660 2516 2518 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08096 2518 2517 2660 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08095 2262 2335 2517 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08094 4478 2338 2262 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08093 4478 2924 2519 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08092 2520 2519 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08091 4478 2436 2519 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08090 2519 2497 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08089 4478 1193 3218 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08088 3218 1189 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08087 3218 1188 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08086 1188 782 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08085 782 716 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08084 4478 721 782 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08083 782 882 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08082 4478 725 782 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08081 4478 715 716 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08080 716 1893 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08079 716 720 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08078 4478 723 721 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08077 721 2934 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08076 721 720 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08075 4478 2488 882 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08074 882 2812 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08073 882 884 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08072 4478 1206 725 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08071 725 2825 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08070 725 724 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08069 1233 1232 1235 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08068 1233 1382 1227 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08067 1227 1225 1233 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08066 1227 1226 1228 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08065 4478 1371 1228 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08064 1235 1396 1233 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08063 1228 1238 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08062 1228 1231 1227 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08061 1237 2229 1238 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08060 4478 1236 1237 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08059 1100 2414 1231 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08058 4478 1101 1100 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08057 1223 1646 1225 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08056 4478 1222 1223 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08055 1397 2410 1396 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08054 4478 1395 1397 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08053 4478 708 1175 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08052 1175 706 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08051 1175 707 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08050 4478 1326 1176 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08049 1176 2809 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08048 1176 1172 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08047 4478 1184 1187 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08046 1189 1187 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08045 4478 1196 1187 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08044 1187 1345 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08043 4478 1357 1196 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08042 1196 2814 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08041 1196 1198 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_08040 1346 1441 1345 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08039 1345 1454 1346 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08038 1346 1343 1344 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08037 1344 1348 1346 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08036 4478 1347 1344 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08035 1344 1451 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08034 1450 1882 1451 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08033 4478 1452 1450 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08032 1342 2175 1343 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08031 4478 1341 1342 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08030 1453 2337 1454 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08029 4478 1452 1453 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_08028 3797 3800 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08027 4478 3808 3800 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08026 3800 3798 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08025 4044 4041 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08024 4478 4329 4044 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08023 4478 4123 4221 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08022 4221 4343 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08021 4221 4122 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08020 4123 4119 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08019 4478 4214 4123 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08018 4478 4341 4346 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08017 4227 4345 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08016 4346 4342 4227 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08015 4338 4333 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08014 4478 4347 4333 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08013 4333 4331 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08012 3913 3914 3912 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_08011 4478 3915 3913 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_08010 4058 3912 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08009 4066 4070 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_08008 4478 4066 3964 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08007 3964 4214 4067 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08006 3682 3916 3803 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_08005 4478 3802 3682 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_08004 4337 3803 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_08003 3916 3915 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_08002 4345 4117 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_08001 4341 4337 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_08000 3917 4058 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07999 3683 3916 3804 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07998 4478 3808 3683 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07997 3963 4067 4064 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07996 4478 4337 3963 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07995 4065 4064 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07994 4478 4058 3961 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07993 3961 4067 3962 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07992 3962 4059 4061 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07991 4122 4061 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07990 3227 3299 4059 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07989 4478 3226 3227 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07988 3906 3908 4053 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07987 4478 3905 3906 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07986 4478 4058 3958 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07985 3958 4338 3957 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07984 3957 4053 4055 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07983 4054 4055 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07982 4478 4044 4210 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07981 4210 4051 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07980 4210 4054 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07979 4226 4338 4340 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07978 4478 4337 4226 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07977 4339 4340 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07976 3909 3911 4056 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07975 4478 3908 3909 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07974 4478 4325 4327 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07973 4327 4332 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07972 4327 4324 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07971 4478 3917 3806 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07970 3684 3808 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07969 3806 3835 3684 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07968 3967 4070 4072 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07967 4478 4071 3967 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07966 4478 3813 3921 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07965 3921 3814 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07964 3921 4068 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07963 4478 4049 4051 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07962 3956 4065 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07961 3956 4320 4049 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07960 4049 4345 3956 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07959 4478 4349 4343 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07958 4228 4346 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07957 4228 4347 4349 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07956 4349 4345 4228 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07955 4478 4336 4332 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07954 4225 4339 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07953 4225 4334 4336 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07952 4336 4345 4225 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07951 4325 4321 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07950 4478 4322 4325 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07949 4478 4058 3959 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07948 3959 4213 3960 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07947 3960 4056 4057 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07946 4324 4057 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07945 3813 3659 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07944 4478 3918 3813 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07943 4478 4337 3966 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07942 3966 4213 3965 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07941 3965 4072 4069 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07940 4068 4069 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07939 4478 3809 3814 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07938 3685 3806 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07937 3685 4334 3809 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07936 3809 3808 3685 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07935 4213 4212 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07934 4478 4320 4212 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07933 4212 4117 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07932 4334 3918 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07931 4320 4322 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07930 4347 4329 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07929 4478 3654 3931 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07928 3931 3654 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07927 4478 3654 3931 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07926 3654 3653 3652 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07925 4478 3804 3654 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07924 3653 3804 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07923 3931 3654 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07922 3654 4214 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07921 4478 3795 4084 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07920 4084 3795 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07919 4478 3795 4084 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07918 3795 3794 3796 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07917 4478 3797 3795 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07916 3794 3797 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07915 4084 3795 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07914 3795 3918 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07913 3792 3790 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07912 4478 3918 3790 4478 tp L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_07911 3904 3903 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07910 4478 4322 3903 4478 tp L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_07909 3907 3910 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07908 4478 4329 3910 4478 tp L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_07907 4218 4214 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07906 4220 4215 4218 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07905 4219 4216 4220 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07904 4217 4216 4223 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07903 4223 4219 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07902 4222 4215 4217 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07901 4216 4118 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07900 4478 4216 4215 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07899 4224 4221 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07898 4478 4224 4222 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07897 4478 4220 4214 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07896 4214 4220 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07895 4219 4217 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07894 4204 4329 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07893 4205 4202 4204 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07892 4208 4203 4205 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07891 4206 4203 4209 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07890 4209 4208 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07889 4207 4202 4206 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07888 4203 4115 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07887 4478 4203 4202 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07886 4211 4210 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07885 4478 4211 4207 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07884 4478 4205 4329 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07883 4329 4205 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07882 4208 4206 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07881 4197 4322 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07880 4311 4319 4197 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07879 4312 4317 4311 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07878 4313 4317 4201 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07877 4201 4312 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07876 4200 4319 4313 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07875 4317 4316 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07874 4478 4317 4319 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07873 4318 4327 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07872 4478 4318 4200 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07871 4478 4311 4322 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07870 4322 4311 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07869 4312 4313 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07868 3919 3918 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07867 3920 3929 3919 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07866 3922 3928 3920 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07865 3925 3928 3924 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07864 3924 3922 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07863 3923 3929 3925 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07862 3928 3926 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07861 4478 3928 3929 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07860 3927 3921 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07859 4478 3927 3923 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07858 4478 3920 3918 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07857 3918 3920 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07856 3922 3925 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07855 3655 3656 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07854 4478 4214 3656 4478 tp L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_07853 3044 3045 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07852 3880 3902 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07851 3269 3209 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07850 3319 3479 3318 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07849 3318 4232 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07848 3317 4107 3319 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07847 4478 3521 3317 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07846 3322 3599 3321 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07845 3321 4107 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07844 3320 4232 3322 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07843 4478 3521 3320 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07842 3254 3073 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07841 3103 3367 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07840 4293 4292 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07839 4269 2786 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07838 4478 3983 3732 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07837 3672 3852 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07836 3732 3729 3672 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07835 4478 3844 3724 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07834 3724 3732 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07833 4478 3733 3724 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07832 3724 3726 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07831 4260 4259 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07830 4164 4163 4165 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07829 4165 4269 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07828 4162 4279 4164 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07827 4478 4161 4162 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07826 3587 3694 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07825 3870 4016 3869 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07824 4478 4167 3870 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07823 3871 3869 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07822 4478 3520 3436 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07821 3436 3515 3521 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07820 3436 3760 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07819 3521 3516 3436 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07818 4478 3760 3515 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07817 3520 3516 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07816 3760 3764 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07815 3764 3766 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07814 4478 3772 3764 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07813 3764 4283 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07812 4478 3771 3764 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07811 4478 4163 3766 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07810 3766 4187 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07809 3766 4196 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07808 3772 3886 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07807 4478 4287 3772 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07806 3771 3774 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07805 4478 4105 3771 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07804 2896 3431 2897 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07803 4478 2916 2896 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07802 2898 2897 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07801 3033 4233 3032 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07800 4478 3031 3033 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07799 3045 3032 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07798 2874 4137 2875 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07797 4478 2873 2874 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07796 2876 2875 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07795 3946 4010 4007 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07794 4478 4186 3946 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07793 4008 4007 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07792 4090 4261 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07791 4478 4269 4090 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07790 4005 4261 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07789 4478 4104 4005 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07788 4240 4241 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07787 4261 4096 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07786 3579 4232 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07785 4478 3584 3580 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07784 3578 3579 3581 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07783 3581 3584 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07782 3581 3580 3578 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07781 4478 4232 3581 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07780 4194 4196 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07779 4478 4198 4195 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07778 4308 4194 4199 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07777 4199 4198 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07776 4199 4195 4308 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07775 4478 4196 4199 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07774 4307 4303 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07773 4478 4308 4309 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07772 4305 4307 4193 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07771 4193 4308 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07770 4193 4309 4305 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07769 4478 4303 4193 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07768 4190 4196 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07767 4478 4198 4189 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07766 4191 4190 4192 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07765 4192 4198 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07764 4192 4189 4191 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07763 4478 4196 4192 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07762 4030 4191 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07761 4478 4032 4037 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07760 4034 4030 3954 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07759 3954 4032 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07758 3954 4037 4034 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07757 4478 4191 3954 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07756 3282 3638 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07755 4478 3635 3283 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07754 3277 3282 3211 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07753 3211 3635 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07752 3211 3283 3277 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07751 4478 3638 3211 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07750 3278 3276 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07749 4478 3277 3275 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07748 3209 3278 3207 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07747 3207 3277 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07746 3207 3275 3209 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07745 4478 3276 3207 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07744 3075 3532 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07743 4478 3075 3076 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07742 3076 3431 3078 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07741 3774 3778 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07740 4478 4298 3778 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07739 3778 3886 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07738 3886 4016 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07737 2882 3503 2883 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07736 4478 2881 2882 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07735 3839 2883 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07734 3840 3698 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07733 4478 4107 3698 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07732 3698 4137 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07731 3072 3781 3071 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07730 4478 3070 3072 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07729 4137 3071 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07728 3785 3787 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07727 4478 4187 3787 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07726 3787 3786 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07725 3681 4039 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07724 3680 3786 3782 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07723 4478 4187 3680 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07722 3782 3785 3681 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07721 3781 3782 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07720 3994 4144 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07719 3941 4024 3998 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07718 4478 4010 3941 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07717 4233 3998 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07716 4028 4029 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07715 4478 4303 4029 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07714 4029 4198 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07713 3953 4039 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07712 3952 4303 4025 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07711 4478 4198 3952 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07710 4025 4028 3953 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07709 4024 4025 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07708 3349 3367 3348 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07707 3346 3344 3349 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07706 3347 3345 3346 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07705 4478 3619 3347 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07704 4478 3348 3506 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07703 3432 3514 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07702 3433 3623 3505 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07701 4478 4269 3433 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07700 3505 3506 3432 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07699 3614 3505 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07698 3345 3343 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07697 4478 3353 3343 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07696 3343 3342 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07695 3357 3355 3356 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07694 4478 3537 3357 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07693 3623 3356 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07692 4262 4258 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07691 2894 3070 2895 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07690 4478 2916 2894 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07689 3499 2895 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07688 2916 2915 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07687 4478 3103 2915 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07686 2915 3786 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07685 3882 3509 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07684 3537 3110 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07683 3514 3510 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07682 4478 3882 3510 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07681 3510 3537 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07680 3619 3710 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07679 4478 3712 3619 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07678 3786 3532 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07677 3354 3509 3353 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07676 4478 3786 3354 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07675 3592 3492 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07674 3583 3255 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07673 4478 3492 3255 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07672 3255 3181 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07671 4478 4269 3179 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07670 3178 3355 3180 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07669 3180 4232 3181 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07668 3179 3514 3178 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07667 3503 3829 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07666 4163 3714 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07665 4302 4301 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07664 4303 4298 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07663 4297 4300 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07662 4478 4298 4300 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07661 4300 4302 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07660 4272 4172 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07659 4478 4105 4172 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07658 4172 4297 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07657 4287 4032 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07656 4285 4289 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07655 4273 4284 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07654 4283 3727 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07653 4177 4283 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07652 4478 4273 4177 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07651 4478 4285 4175 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07650 4175 4283 4176 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07649 4176 4284 4286 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07648 4295 4286 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07647 4280 4015 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07646 4478 4032 4015 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07645 4015 4273 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07644 4279 4281 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07643 4478 4280 4281 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07642 4281 4290 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07641 4186 4185 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07640 4478 4273 4185 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07639 4185 4303 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07638 4167 4104 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07637 3949 4301 4011 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07636 3948 4167 3949 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07635 3947 4186 3948 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07634 4478 4163 3947 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07633 4478 4011 4161 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07632 3951 4196 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07631 3950 4287 4018 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07630 4478 4187 3950 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07629 4018 4020 3951 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07628 4146 4018 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07627 4020 4022 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07626 4478 4187 4022 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07625 4022 4287 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07624 4149 4146 4148 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07623 4478 4272 4149 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07622 3667 3983 3696 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07621 4478 3690 3667 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07620 3694 3696 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07619 3439 4196 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07618 3438 3537 3525 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07617 4478 4198 3438 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07616 3525 3531 3439 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07615 3526 3525 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07614 3531 3529 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07613 4478 3537 3529 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07612 3529 4198 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07611 3325 3331 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07610 3596 3594 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07609 4478 3727 3597 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07608 3599 3596 3598 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07607 3598 3727 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07606 3598 3597 3599 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07605 4478 3594 3598 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07604 4478 4296 4183 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07603 4182 4179 4183 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07602 4183 4180 4182 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07601 4478 4294 4184 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07600 4181 4295 4296 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07599 4184 4293 4181 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07598 4010 4013 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07597 4478 4105 4013 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07596 4013 4280 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07595 2919 2918 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07594 4478 3110 2918 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07593 2918 3103 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07592 3070 2800 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07591 4105 4038 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07590 3846 3502 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07589 4243 2886 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07588 4107 4232 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07587 4187 4198 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07586 3636 3638 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07585 3983 3991 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07584 4039 4196 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07583 3637 3635 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07582 4147 4272 4259 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07581 4478 4285 4147 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07580 4153 4261 4278 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07579 4478 4262 4153 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07578 3310 3171 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07577 4478 4107 3310 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07576 4140 4252 4258 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07575 4478 4253 4140 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07574 3942 3999 4104 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07573 4478 4102 3942 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07572 4136 4261 4241 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07571 4478 4253 4136 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07570 4478 3705 3668 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07569 3668 3709 4096 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07568 3668 3710 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07567 4096 3712 3668 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07566 4478 3710 3709 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07565 3705 3712 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07564 3239 4233 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07563 4478 4269 3239 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07562 2868 2867 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07561 4478 4269 2867 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07560 2867 4137 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07559 4478 3899 3901 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07558 3901 3900 3902 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07557 3901 4198 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07556 3902 4196 3901 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07555 4478 4198 3900 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07554 3899 4196 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07553 4478 3077 3074 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07552 3073 4105 3074 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07551 3074 3078 3073 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07550 4016 4163 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07549 4478 4302 4016 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07548 3431 3882 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07547 4478 3503 3431 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07546 3582 4148 3584 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07545 4478 3594 3582 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07544 3492 3353 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07543 4478 4105 3492 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07542 2893 4269 3331 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07541 4478 3619 2893 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07540 3744 3747 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07539 4478 4283 3747 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07538 3747 3745 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07537 3863 4280 3862 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07536 4478 3871 3863 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07535 3864 3862 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07534 3675 4269 3741 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07533 4478 4280 3675 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07532 3742 3741 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07531 3193 3189 3262 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07530 3193 3190 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07529 4478 3625 3193 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07528 3262 3846 3193 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07527 3188 3262 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07526 4478 3082 3189 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07525 3189 3098 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07524 3189 3083 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07523 4478 3077 3079 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07522 3079 3091 3080 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07521 3080 3078 3081 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07520 3083 3081 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07519 4478 4269 3082 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07518 3082 2890 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07517 3082 3983 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07516 4478 2885 2887 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07515 2887 2888 2890 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07514 2887 4232 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07513 2890 2886 2887 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07512 4478 4232 2888 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07511 2885 2886 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07510 4478 3096 3101 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07509 3101 3774 3100 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07508 3100 4243 3102 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07507 3098 3102 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07506 4478 4111 3625 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07505 3625 3630 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07504 3625 3624 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07503 4478 3633 3624 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07502 3624 3623 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07501 3624 3626 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07500 4478 4243 4111 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07499 4111 4113 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07498 4478 4179 4113 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07497 4478 3991 3630 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07496 3631 3634 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07495 3630 3629 3631 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07494 3632 3633 3634 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07493 4478 4102 3632 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07492 4478 3633 3628 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07491 3629 3628 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07490 4478 3627 3628 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07489 3628 4102 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07488 4098 4232 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07487 4478 4233 4098 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07486 4145 4163 4144 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07485 4478 4143 4145 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07484 3711 3710 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07483 4478 3711 3670 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07482 3670 3712 3714 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07481 2800 2919 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07480 4478 4105 2800 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07479 3669 3712 3829 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07478 4478 3710 3669 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07477 4178 4287 4179 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07476 4478 4177 4178 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07475 4292 4290 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07474 4478 4297 4292 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07473 4298 3638 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07472 4478 3637 4298 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07471 4289 4287 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07470 4478 4302 4289 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07469 4188 4187 4301 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07468 4478 4196 4188 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07467 4032 3635 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07466 4478 3636 4032 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07465 3955 4039 4284 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07464 4478 4198 3955 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07463 3601 3712 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07462 4478 3601 3600 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07461 3600 3710 3727 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07460 3355 3619 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07459 4478 3103 3355 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07458 3532 3636 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07457 4478 3637 3532 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07456 3437 4196 3509 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07455 4478 4198 3437 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07454 3110 3638 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07453 4478 3635 3110 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07452 3367 3366 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07451 4478 4196 3366 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07450 3366 4198 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07449 4478 3835 2787 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07448 2788 3911 2789 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07447 2789 3226 2790 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07446 2787 3905 2788 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07445 3658 3657 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07444 4478 3835 3657 4478 tp L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_07443 3867 4010 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07442 3866 4182 3868 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07441 4478 4107 3866 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07440 3868 4161 3867 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07439 3865 3868 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07438 3674 4243 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07437 3673 4269 3736 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07436 4478 3735 3673 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07435 3736 3865 3674 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07434 3733 3736 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07433 3620 3619 3621 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07432 4478 4167 3620 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07431 3615 4107 3616 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07430 4478 3614 3615 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07429 4478 3617 3729 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07428 3617 4243 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07427 4478 3616 3618 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07426 3618 3621 3617 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07425 3943 4182 4001 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07424 4478 4102 3943 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07423 4155 4283 4263 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07422 4478 4262 4155 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07421 4478 3854 3852 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07420 3854 3850 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07419 4478 4263 3853 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07418 3853 4001 3854 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07417 4478 4144 4141 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07416 4142 4141 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07415 4478 4101 4141 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07414 4141 4098 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07413 4478 3850 3841 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07412 3842 3839 3843 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07411 3841 3840 3842 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07410 4478 3991 3844 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07409 3845 3843 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07408 3844 4142 3845 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07407 4478 4262 3427 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07406 3428 3499 3429 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07405 3429 3509 3606 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07404 3427 3503 3428 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07403 3609 3614 3608 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07402 4478 4102 3609 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07401 4478 4243 3726 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07400 3607 3608 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07399 3726 3606 3607 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07398 4478 4294 4159 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07397 4160 4295 4264 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07396 4159 4272 4160 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07395 4478 4269 4156 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07394 4158 4177 4157 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07393 4156 4260 4158 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07392 4478 4154 4152 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07391 4154 4102 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07390 4478 4157 4103 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07389 4103 4264 4154 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07388 4478 4243 4150 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07387 4151 4164 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07386 4150 4152 4151 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07385 3486 3326 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07384 4478 3325 3326 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07383 3326 3327 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07382 4478 3526 3418 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07381 3420 3592 3489 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07380 3418 4269 3420 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07379 4478 3487 3488 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07378 3487 3486 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07377 4478 3489 3417 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07376 3417 4107 3487 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07375 3410 4148 3466 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07374 4478 4232 3410 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07373 3468 3466 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07372 4478 3468 3467 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07371 3470 3467 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07370 4478 4243 3467 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07369 3467 3599 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07368 4478 3983 3701 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07367 3413 3470 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07366 3701 3488 3413 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07365 3593 3592 3595 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07364 4478 3594 3593 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07363 4478 4232 3591 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07362 3591 3585 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07361 4478 3584 3585 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07360 3589 3591 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07359 4478 3587 3589 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07358 3589 3714 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07357 3589 3583 3590 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07356 3590 3829 3588 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07355 3700 3586 3589 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07354 3588 3595 3700 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07353 4478 3701 3716 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07352 3716 4150 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07351 3716 3700 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07350 3671 3716 3720 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07349 3671 3846 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07348 4478 3724 3671 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07347 3720 3717 3671 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07346 3715 3720 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07345 2869 2868 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07344 3038 3239 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07343 3677 3754 3752 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07342 4478 3749 3678 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07341 3676 3846 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07340 3752 3872 3676 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07339 3678 3748 3677 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07338 3679 3887 3678 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07337 3752 4243 3679 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07336 3905 3752 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07335 3754 4243 4478 4478 tp L=0.32U W=1.9U AS=1.425P AD=1.425P PS=5.3U PD=5.3U 
Mtr_07334 4478 3846 3749 4478 tp L=0.32U W=1.9U AS=1.425P AD=1.425P PS=5.3U PD=5.3U 
Mtr_07333 3878 3875 3877 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07332 4478 3874 3879 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07331 3873 4243 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07330 3877 3881 3873 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07329 3879 3896 3878 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07328 3876 3880 3879 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07327 3877 4269 3876 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07326 3872 3877 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07325 3875 4269 4478 4478 tp L=0.32U W=1.9U AS=1.425P AD=1.425P PS=5.3U PD=5.3U 
Mtr_07324 4478 4243 3874 4478 tp L=0.32U W=1.9U AS=1.425P AD=1.425P PS=5.3U PD=5.3U 
Mtr_07323 3885 3902 3883 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07322 3885 4269 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07321 4478 3882 3885 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07320 3883 3884 3885 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07319 3881 3883 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07318 3896 4034 3898 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07317 3898 4105 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07316 3897 3895 3896 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07315 4478 4305 3897 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07314 3361 3363 3360 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07313 4478 3358 3364 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07312 3359 4269 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07311 3360 3367 3359 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07310 3364 3370 3361 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07309 3365 3538 3364 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07308 3360 3362 3365 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07307 3748 3360 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07306 3363 3362 4478 4478 tp L=0.32U W=1.9U AS=1.425P AD=1.425P PS=5.3U PD=5.3U 
Mtr_07305 4478 4269 3358 4478 tp L=0.32U W=1.9U AS=1.425P AD=1.425P PS=5.3U PD=5.3U 
Mtr_07304 3368 3372 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07303 4478 3532 3369 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07302 3370 3368 3371 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07301 3371 3532 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07300 3371 3369 3370 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07299 4478 3372 3371 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07298 3373 4196 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07297 4478 4198 3375 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07296 3372 3373 3374 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07295 3374 4198 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07294 3374 3375 3372 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07293 4478 4196 3374 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07292 3534 3537 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07291 4478 3548 3535 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07290 3538 3534 3441 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07289 3441 3548 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07288 3441 3535 3538 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07287 4478 3537 3441 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07286 3542 4196 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07285 4478 4198 3543 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07284 3548 3542 3443 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07283 3443 4198 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07282 3443 3543 3548 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07281 4478 4196 3443 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07280 3892 3893 3891 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07279 4478 3888 3894 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07278 3890 4269 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07277 3891 4284 3890 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07276 3894 4034 3892 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07275 3889 4305 3894 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07274 3891 4105 3889 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07273 3887 3891 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07272 3893 4105 4478 4478 tp L=0.35U W=1.9U AS=1.463P AD=1.463P PS=5.35U PD=5.35U 
Mtr_07271 4478 4269 3888 4478 tp L=0.35U W=1.9U AS=1.463P AD=1.463P PS=5.35U PD=5.35U 
Mtr_07270 3090 3087 3089 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07269 4478 3086 3095 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07268 3088 3084 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07267 3089 3194 3088 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07266 3095 3085 3090 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07265 3093 3109 3095 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07264 3089 3091 3093 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07263 3226 3089 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07262 3087 3091 4478 4478 tp L=0.32U W=1.9U AS=1.425P AD=1.425P PS=5.3U PD=5.3U 
Mtr_07261 4478 3084 3086 4478 tp L=0.32U W=1.9U AS=1.425P AD=1.425P PS=5.3U PD=5.3U 
Mtr_07260 3094 3201 3197 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07259 4478 3195 3099 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07258 3092 4243 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07257 3197 3200 3092 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07256 3099 3209 3094 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07255 3097 3537 3099 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07254 3197 4269 3097 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07253 3194 3197 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07252 3201 4269 4478 4478 tp L=0.32U W=1.9U AS=1.425P AD=1.425P PS=5.3U PD=5.3U 
Mtr_07251 4478 4243 3195 4478 tp L=0.32U W=1.9U AS=1.425P AD=1.425P PS=5.3U PD=5.3U 
Mtr_07250 4478 3270 3200 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07249 3204 4287 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07248 3268 3272 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07247 3203 3272 3270 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07246 3270 3268 3204 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07245 4478 3269 3203 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07244 3085 2944 2921 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07243 2921 4269 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07242 2920 2926 3085 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07241 4478 3786 2920 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07240 2943 3635 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07239 4478 3638 2946 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07238 2944 2943 2945 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07237 2945 3638 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07236 2945 2946 2944 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07235 4478 3635 2945 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07234 4478 3104 3108 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07233 3108 3107 3109 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07232 3108 3106 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07231 3109 3105 3108 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07230 4478 3106 3107 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07229 3104 3105 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07228 2938 3638 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07227 4478 3635 2941 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07226 3106 2938 2939 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07225 2939 3635 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07224 2939 2941 3106 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07223 4478 3638 2939 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07222 2927 2926 2928 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07221 4478 2925 2927 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07220 3105 2928 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07219 3061 3057 3059 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07218 4478 3056 3060 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07217 3054 3055 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07216 3059 3065 3054 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07215 3060 3158 3061 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07214 3058 3165 3060 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07213 3059 3991 3058 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07212 4397 3059 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07211 3057 3991 4478 4478 tp L=0.32U W=1.9U AS=1.425P AD=1.425P PS=5.3U PD=5.3U 
Mtr_07210 4478 3055 3056 4478 tp L=0.32U W=1.9U AS=1.425P AD=1.425P PS=5.3U PD=5.3U 
Mtr_07209 3065 3069 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07208 4478 3064 3067 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07207 3067 3991 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07206 3067 3855 3068 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07205 3068 3091 3067 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07204 3069 4243 3068 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07203 3068 3066 3069 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07202 3064 3052 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07201 4478 3053 3064 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07200 4478 3994 3052 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07199 3052 3048 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07198 3052 3049 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07197 3048 4232 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07196 4478 3045 3048 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07195 4478 3839 3053 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07194 3053 2878 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07193 3053 4243 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07192 2878 2876 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07191 4478 4107 2878 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07190 4478 3861 3855 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07189 3855 3858 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07188 3855 4283 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07187 3860 3871 3859 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07186 4478 4008 3860 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07185 3861 3859 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07184 3857 4269 3856 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07183 4478 4010 3857 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07182 3858 3856 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07181 4478 2792 3066 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07180 3066 2798 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07179 3066 3619 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07178 4478 3253 2793 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07177 2793 3070 2791 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07176 2791 2898 2794 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07175 2792 2794 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07174 2798 2799 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07173 4478 2800 2798 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07172 4478 3247 3158 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07171 3157 3164 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07170 3157 3319 3247 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07169 3247 4243 3157 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07168 4478 3475 3414 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07167 3414 3476 3479 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07166 3414 3714 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07165 3479 3477 3414 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07164 4478 3714 3476 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07163 3475 3477 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07162 4478 3583 3163 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07161 3162 3161 3164 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07160 3163 4243 3162 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07159 4478 3073 3063 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07158 3161 3503 3063 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07157 3063 3062 3161 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07156 3165 3169 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07155 3167 3177 3166 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07154 3167 4243 4478 4478 tp L=0.32U W=4.05U AS=3.0375P AD=3.0375P PS=9.6U PD=9.6U 
Mtr_07153 4478 3322 3167 4478 tp L=0.32U W=4.05U AS=3.0375P AD=3.0375P PS=9.6U PD=9.6U 
Mtr_07152 3166 3174 3169 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07151 3169 3172 3167 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07150 4478 3325 3174 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07149 3174 3254 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07148 3174 4167 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07147 4478 4269 2795 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07146 2796 2900 2797 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07145 2797 4107 3177 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07144 2795 2898 2796 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07143 2900 2901 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07142 4478 2919 2901 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07141 2901 2925 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07140 4478 3498 3493 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07139 3421 3495 3498 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07138 3422 3847 3421 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07137 3423 3983 3422 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07136 3423 3496 4478 4478 tp L=0.35U W=3.05U AS=2.3485P AD=2.3485P PS=7.65U PD=7.65U 
Mtr_07135 4478 3502 3423 4478 tp L=0.35U W=3.05U AS=2.3485P AD=2.3485P PS=7.65U PD=7.65U 
Mtr_07134 3423 3603 4478 4478 tp L=0.35U W=3.05U AS=2.3485P AD=2.3485P PS=7.65U PD=7.65U 
Mtr_07133 3498 3613 3423 4478 tp L=0.35U W=3.32U AS=2.5564P AD=2.5564P PS=8.2U PD=8.2U 
Mtr_07132 3496 3622 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07131 4478 3507 3496 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07130 4478 4163 3622 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07129 3622 4174 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07128 3622 4243 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07127 4478 4177 4109 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07126 4109 4297 4108 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07125 4108 4107 4173 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07124 4174 4173 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07123 4478 3352 3507 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07122 3507 3258 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07121 3507 3260 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07120 3187 3353 3261 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07119 4478 3272 3187 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07118 3260 3261 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07117 3352 3351 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07116 4478 3503 3351 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07115 3351 3350 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07114 4478 3310 3183 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07113 3183 3353 3184 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07112 3184 3355 3257 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07111 3258 3257 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07110 4478 3602 3603 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07109 3603 3604 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07108 3603 3983 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07107 4478 3327 3602 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07106 3328 3329 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07105 3602 3331 3328 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07104 4478 4107 3330 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07103 3329 3781 3330 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07102 3330 3344 3329 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07101 4478 4243 3604 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07100 3605 3851 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07099 3604 3727 3605 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07098 3848 4024 3851 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07097 4478 4102 3848 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07096 4478 3482 3416 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07095 3495 3481 3416 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07094 3416 3839 3495 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07093 4478 3323 3481 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07092 3324 4232 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07091 3324 4269 3323 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07090 3323 3526 3324 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07089 4478 4243 3849 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07088 3847 3996 3849 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07087 3849 3994 3847 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07086 4478 3997 3996 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07085 3940 4252 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07084 3940 4269 3997 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07083 3997 4146 3940 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07082 4478 3610 3612 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07081 3613 3611 3612 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07080 3612 3740 3613 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07079 4478 2907 3611 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07078 3611 2905 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07077 3611 2913 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07076 2913 2912 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07075 4478 4243 2912 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07074 2912 3619 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07073 2909 4269 2910 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07072 4478 2919 2909 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07071 2907 2910 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07070 4478 3253 2902 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07069 2902 2919 2903 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07068 2903 3431 2904 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07067 2905 2904 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07066 4478 3864 3740 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07065 3740 3742 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07064 3740 3744 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07063 3835 3837 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07062 3838 3833 3834 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07061 3838 3846 4478 4478 tp L=0.35U W=4.05U AS=3.1185P AD=3.1185P PS=9.65U PD=9.65U 
Mtr_07060 4478 3981 3838 4478 tp L=0.35U W=4.05U AS=3.1185P AD=3.1185P PS=9.65U PD=9.65U 
Mtr_07059 3834 4246 3837 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07058 3837 3836 3838 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07057 3981 3988 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07056 3936 4092 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07055 4478 3983 3936 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07054 3936 3991 3937 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07053 3988 3990 3938 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07052 3937 3982 3936 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07051 3937 4243 3938 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07050 3938 3986 3937 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07049 3938 4265 3988 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07048 4092 4238 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07047 4478 4135 4092 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07046 4478 4241 4238 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07045 4238 4236 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07044 4238 4235 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07043 4133 4233 4234 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07042 4478 4232 4133 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07041 4236 4234 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07040 4478 4088 4089 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07039 4089 4090 4091 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07038 4091 4139 4134 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07037 4135 4134 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07036 4138 4252 4139 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07035 4478 4137 4138 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07034 3982 3973 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07033 4478 4132 3982 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_07032 4478 3840 3818 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07031 3818 3819 3817 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07030 3817 4240 3820 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07029 3973 3820 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07028 4478 4243 4086 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07027 4086 4090 4085 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07026 4085 4094 4131 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07025 4132 4131 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07024 4094 4098 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07023 4478 3331 3332 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07022 3332 3341 3333 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07021 3333 3336 3334 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07020 3986 3334 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_07019 4478 3345 3338 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07018 3339 3514 3340 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07017 3340 3367 3341 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07016 3338 4005 3339 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07015 4478 3499 3335 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07014 3337 4003 3336 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07013 3335 3509 3337 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07012 4003 4278 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07011 4478 4275 4265 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07010 4265 4266 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07009 4265 4270 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07008 4166 4269 4271 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07007 4478 4283 4166 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_07006 4270 4271 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_07005 4478 4292 4275 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07004 4275 4273 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07003 4478 4289 4275 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07002 4275 4278 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_07001 4478 4008 3945 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_07000 3945 4005 3944 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06999 3944 4301 4006 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06998 4266 4006 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06997 4246 4245 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06996 4478 4243 4245 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06995 4245 4250 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06994 4478 4256 4250 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06993 4250 4248 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06992 4250 4247 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06991 4247 4253 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06990 4478 4261 4247 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06989 4478 4259 4256 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06988 4256 4261 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06987 4478 4258 4256 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06986 4256 4273 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06985 4248 4096 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06984 4478 4169 4248 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06983 4478 4186 4168 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06982 4171 4167 4170 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06981 4170 4279 4169 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06980 4168 4301 4171 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06979 4478 3972 3833 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06978 3833 3824 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06977 3833 3823 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06976 4478 3694 3665 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_06975 3665 4240 3666 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_06974 3666 3691 3692 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_06973 3823 3692 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06972 3691 3689 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06971 4478 4148 3689 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06970 3689 4232 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06969 4478 3980 3972 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06968 3934 4232 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06967 3972 3977 3934 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06966 3977 3979 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06965 4478 4269 3979 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06964 3979 4148 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06963 3978 4261 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06962 4478 3978 3935 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06961 3935 3993 3980 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06960 3939 3990 3992 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06959 4478 3991 3939 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06958 3993 3992 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06957 4478 3827 3824 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06956 3826 4243 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06955 3826 3832 3827 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06954 3827 3825 3826 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06953 3831 3829 3830 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_06952 4478 3828 3831 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_06951 3832 3830 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06950 3821 4269 3822 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_06949 4478 4261 3821 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_06948 3825 3822 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06947 3046 3156 3150 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06946 4478 3149 3050 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06945 3047 3846 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06944 3150 3303 3047 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06943 3050 3152 3046 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06942 3051 3153 3050 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06941 3150 3991 3051 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06940 3911 3150 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06939 3156 3991 4478 4478 tp L=0.35U W=1.9U AS=1.463P AD=1.463P PS=5.35U PD=5.35U 
Mtr_06938 4478 3846 3149 4478 tp L=0.35U W=1.9U AS=1.463P AD=1.463P PS=5.35U PD=5.35U 
Mtr_06937 3309 3305 3308 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06936 4478 3304 3306 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06935 3302 3983 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06934 3308 3312 3302 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06933 3306 3578 3309 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06932 3307 3460 3306 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06931 3308 4243 3307 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06930 3303 3308 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06929 3305 4243 4478 4478 tp L=0.35U W=1.9U AS=1.463P AD=1.463P PS=5.35U PD=5.35U 
Mtr_06928 4478 3983 3304 4478 tp L=0.35U W=1.9U AS=1.463P AD=1.463P PS=5.35U PD=5.35U 
Mtr_06927 4478 3316 3312 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06926 3311 3310 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06925 3314 3327 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06924 3315 3327 3316 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06923 3316 3314 3311 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06922 4478 3313 3315 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06921 3313 3578 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_06920 3458 3463 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06919 4478 4232 3459 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06918 3460 3458 3409 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06917 3409 4232 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06916 3409 3459 3460 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06915 4478 3463 3409 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06914 3146 3145 3243 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06913 3146 3144 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06912 4478 3142 3146 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06911 3243 4243 3146 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06910 3152 3243 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06909 2862 4232 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06908 4478 2868 2865 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06907 3145 2862 2863 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06906 2863 2868 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06905 2863 2865 3145 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06904 4478 4232 2863 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06903 3236 4232 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06902 4478 3239 3237 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06901 3142 3236 3139 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06900 3139 3239 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06899 3139 3237 3142 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06898 4478 4232 3139 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06897 3043 3037 3042 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06896 4478 3039 3040 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06895 3036 3035 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06894 3042 3034 3036 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06893 3040 3038 3043 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06892 3041 3044 3040 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06891 3042 4107 3041 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06890 3153 3042 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06889 3037 4107 4478 4478 tp L=0.35U W=1.9U AS=1.463P AD=1.463P PS=5.35U PD=5.35U 
Mtr_06888 4478 3035 3039 4478 tp L=0.35U W=1.9U AS=1.463P AD=1.463P PS=5.35U PD=5.35U 
Mtr_06887 3034 2869 2871 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06886 2871 4107 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06885 2870 4232 3034 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06884 4478 2876 2870 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06883 3393 3390 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06882 3392 3393 3391 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06881 4478 3394 3392 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06880 2951 3397 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06879 2965 3390 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06878 2967 2965 2968 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06877 4478 2966 2967 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06876 2966 2963 2962 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06875 2962 3226 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06874 2961 3221 2966 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06873 4478 3397 2961 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06872 2963 3397 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06871 3131 3130 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06870 4478 3390 3130 4478 tp L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_06869 2974 2973 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06868 4478 2971 2973 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06867 2973 2970 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06866 3449 3570 4352 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06865 4478 3569 3449 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06864 3390 3234 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_06863 3570 3568 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06862 4478 3398 3400 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06861 3400 3399 3402 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06860 3402 3404 3401 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06859 3397 3401 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06858 3404 3403 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_06857 2957 2951 2949 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06856 2949 3905 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06855 2948 3380 2957 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06854 4478 3397 2948 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06853 2956 3390 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06852 2958 2956 2959 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06851 4478 2957 2958 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06850 2954 3397 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_06849 3127 2954 2953 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06848 2953 3911 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06847 2952 3218 3127 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06846 4478 3397 2952 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06845 3126 3390 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06844 3129 3126 3128 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06843 4478 3127 3129 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06842 3562 3560 4478 4478 tp L=0.35U W=4.2U AS=3.234P AD=3.234P PS=9.95U PD=9.95U 
Mtr_06841 3561 3567 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06840 4478 3570 3563 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06839 3563 3561 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06838 4478 3562 3563 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06837 3563 3569 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06836 3396 3397 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06835 4478 3563 3394 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06834 3395 3396 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06833 3394 3835 3395 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06832 3710 3646 3649 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06831 3649 3799 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06830 3648 3647 3710 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06829 4478 3651 3648 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06828 3219 3447 3288 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06827 3219 4458 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06826 4478 3220 3219 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06825 3288 3218 3219 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06824 4102 3288 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06823 4478 3382 4198 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06822 3381 3386 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06821 3381 3447 3382 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06820 3382 3380 3381 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06819 3222 3447 3292 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06818 3222 4470 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06817 4478 3225 3222 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06816 3292 3221 3222 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06815 3638 3292 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06814 4478 3639 3712 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06813 3712 3645 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06812 3712 3641 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06811 4478 3792 3641 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06810 3641 3640 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06809 4478 3643 3640 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06808 4478 3114 3991 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06807 3991 3112 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06806 3991 3113 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06805 3558 3560 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06804 4478 3558 3448 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06803 3448 3559 3650 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06802 3446 3647 3447 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06801 4478 3559 3446 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06800 4478 3389 3119 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06799 3119 3122 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06798 3119 3118 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06797 3120 3221 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06796 4478 3553 3120 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06795 4478 3123 3635 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06794 3635 3119 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06793 3635 3120 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06792 4478 3907 3642 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06791 3642 3644 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06790 4478 3643 3644 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06789 3379 3380 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06788 4478 3553 3379 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06787 4478 3642 4196 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06786 4196 3378 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06785 4196 3379 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06784 3799 4452 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06783 3651 3650 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06782 3220 3646 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06781 3225 3646 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06780 3555 3286 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06779 3554 3559 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06778 3389 3647 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06777 3553 3550 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06776 4478 3554 3550 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06775 3550 3647 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06774 3385 3553 3384 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06773 4478 3383 3385 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06772 3643 3384 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06771 4478 3445 3646 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06770 3646 3388 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06769 4478 3389 3388 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06768 4478 3445 3387 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06767 3386 3387 4478 4478 tp L=0.35U W=5.62U AS=4.3274P AD=4.3274P PS=12.8U PD=12.8U 
Mtr_06766 4478 4464 3387 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06765 3387 3647 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06764 4478 3286 3639 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06763 3639 3389 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06762 3639 3289 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06761 3116 3643 3115 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06760 4478 3793 3116 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06759 3114 3115 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_06758 4478 3389 3112 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06757 3112 3117 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06756 3112 3111 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06755 4478 3555 3122 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06754 3122 3121 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06753 4478 3655 3121 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06752 3445 3554 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06751 4478 3555 3445 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06750 4478 3553 3124 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06749 3124 3125 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06748 4478 3221 3125 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06747 4478 3555 3123 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06746 3123 3124 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06745 3123 3655 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06744 4478 3376 3378 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06743 3378 3389 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06742 3378 3377 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06741 3645 3647 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06740 4478 3650 3645 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06739 3113 3218 4478 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06738 4478 3553 3113 4478 tp L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_06737 3793 3904 4478 4478 tp L=0.32U W=4.2U AS=3.15P AD=3.15P PS=9.9U PD=9.9U 
Mtr_06736 3117 3793 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_06735 4478 3555 3117 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.p17d 4478 4468 4469 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.p14d 4535 4531 4545 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_d0.p18f 4478 4469 4470 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d0.p18d 4478 4469 4470 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d0.p2 4467 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.p17a 4469 4468 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.p0 4478 4540 4466 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.p4b 4478 4467 4494 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.p14b 4535 4531 4545 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_d0.p16 4468 4469 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_d0.p17b 4478 4468 4469 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.p4a 4494 4467 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.p18a 4470 4469 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d0.p18e 4470 4469 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d0.p3 4465 4466 4467 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.p7c 4533 4493 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d0.p5a 4493 4465 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.p7b 4535 4493 4533 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d0.p7a 4533 4493 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d0.p10 4535 4531 4530 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d0.p13 4530 4545 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d0.p6c 4535 4494 4532 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d0.p6b 4532 4494 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d0.p6a 4535 4494 4532 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d0.p8c 4532 4545 4531 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d0.p14c 4545 4531 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_d0.p8b 4531 4545 4532 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d0.p18b 4478 4469 4470 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d0.p17c 4469 4468 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.p8a 4532 4545 4531 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d0.p9 4531 4535 4545 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d0.p12 4545 4535 4530 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d0.p5b 4478 4465 4493 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.p1 4478 4540 4467 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.p14a 4545 4531 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_d0.p11 4545 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_d0.p18c 4470 4469 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d1.p17d 4478 4462 4463 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.p14d 4535 4527 4544 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_d1.p18f 4478 4463 4464 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d1.p18d 4478 4463 4464 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d1.p2 4461 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.p17a 4463 4462 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.p0 4478 4540 4460 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.p4b 4478 4461 4492 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.p14b 4535 4527 4544 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_d1.p16 4462 4463 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_d1.p17b 4478 4462 4463 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.p4a 4492 4461 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.p18a 4464 4463 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d1.p18e 4464 4463 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d1.p3 4459 4460 4461 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.p7c 4528 4491 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d1.p5a 4491 4459 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.p7b 4535 4491 4528 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d1.p7a 4528 4491 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d1.p10 4535 4527 4525 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d1.p13 4525 4544 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d1.p6c 4535 4492 4526 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d1.p6b 4526 4492 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d1.p6a 4535 4492 4526 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d1.p8c 4526 4544 4527 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d1.p14c 4544 4527 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_d1.p8b 4527 4544 4526 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d1.p18b 4478 4463 4464 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d1.p17c 4463 4462 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.p8a 4526 4544 4527 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d1.p9 4527 4535 4544 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d1.p12 4544 4535 4525 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d1.p5b 4478 4459 4491 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.p1 4478 4540 4461 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.p14a 4544 4527 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_d1.p11 4544 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_d1.p18c 4464 4463 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i7.p17d 4478 60 61 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.p14d 4535 6 9 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i7.p18f 4478 61 123 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i7.p18d 4478 61 123 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i7.p2 56 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.p17a 61 60 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.p0 4478 4540 55 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.p4b 4478 56 58 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.p14b 4535 6 9 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i7.p16 60 61 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_i7.p17b 4478 60 61 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.p4a 58 56 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.p18a 123 61 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i7.p18e 123 61 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i7.p3 57 55 56 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.p7c 10 54 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i7.p5a 54 57 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.p7b 4535 54 10 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i7.p7a 10 54 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i7.p10 4535 6 7 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i7.p13 7 9 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i7.p6c 4535 58 8 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i7.p6b 8 58 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i7.p6a 4535 58 8 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i7.p8c 8 9 6 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i7.p14c 9 6 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i7.p8b 6 9 8 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i7.p18b 4478 61 123 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i7.p17c 61 60 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.p8a 8 9 6 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i7.p9 6 4535 9 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i7.p12 9 4535 7 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i7.p5b 4478 57 54 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.p1 4478 4540 56 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.p14a 9 6 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_i7.p11 9 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_i7.p18c 123 61 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_ovr.p17a 1662 1663 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.p18d 4478 1662 1550 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_ovr.p14d 4535 1942 1828 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_ovr.p18f 4478 1662 1550 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_ovr.p18c 1550 1662 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_ovr.p17d 4478 1663 1662 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.p11 1828 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_ovr.p14a 1828 1942 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_ovr.p1 4478 3715 1829 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.p12 1828 4535 1943 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ovr.p9 1942 4535 1828 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ovr.p5b 4478 1830 1832 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.p8a 1693 1828 1942 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ovr.p8b 1942 1828 1693 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ovr.p8c 1693 1828 1942 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ovr.p14c 1828 1942 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_ovr.p6a 4535 1695 1693 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ovr.p18b 4478 1662 1550 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_ovr.p6b 1693 1695 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ovr.p6c 4535 1695 1693 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ovr.p17c 1662 1663 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.p13 1943 1828 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ovr.p10 4535 1942 1943 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ovr.p7a 1694 1832 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ovr.p7b 4535 1832 1694 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ovr.p7c 1694 1832 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ovr.p3 1830 1831 1829 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.p5a 1832 1830 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.p4a 1695 1829 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.p18a 1550 1662 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_ovr.p18e 1550 1662 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_ovr.p17b 4478 1663 1662 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.p16 1663 1662 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_ovr.p14b 4535 1942 1828 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_ovr.p4b 4478 1829 1695 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.p0 4478 4478 1831 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.p2 1829 4478 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.p17d 4478 4441 4442 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.p18c 4443 4442 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y0.p18f 4478 4442 4443 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y0.p14d 4535 4511 4539 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_y0.p18d 4478 4442 4443 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y0.p2 4440 4437 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.p17a 4442 4441 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.p4b 4478 4440 4486 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.p0 4478 4437 4439 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.p16 4441 4442 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_y0.p14b 4535 4511 4539 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_y0.p17b 4478 4441 4442 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.p4a 4486 4440 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.p7c 4513 4485 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y0.p18e 4443 4442 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y0.p7b 4535 4485 4513 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y0.p18a 4443 4442 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y0.p7a 4513 4485 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y0.p10 4535 4511 4510 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y0.p3 4438 4439 4440 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.p13 4510 4539 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y0.p5a 4485 4438 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.p6c 4535 4486 4512 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y0.p6b 4512 4486 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y0.p6a 4535 4486 4512 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y0.p8c 4512 4539 4511 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y0.p8b 4511 4539 4512 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y0.p17c 4442 4441 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.p8a 4512 4539 4511 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y0.p9 4511 4535 4539 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y0.p12 4539 4535 4510 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y0.p14c 4539 4511 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_y0.p18b 4478 4442 4443 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y0.p1 4478 4436 4440 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.p5b 4478 4438 4485 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.p14a 4539 4511 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_y0.p11 4539 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_b0.p17d 4478 1278 1398 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.p14d 4535 1242 1402 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_b0.p18f 4478 1398 1399 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b0.p18d 4478 1398 1399 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b0.p2 1104 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.p17a 1398 1278 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.p0 4478 4540 994 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.p4b 4478 1104 1240 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.p14b 4535 1242 1402 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_b0.p16 1278 1398 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_b0.p17b 4478 1278 1398 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.p4a 1240 1104 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.p18a 1399 1398 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b0.p18e 1399 1398 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b0.p3 993 994 1104 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.p7c 1400 1239 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b0.p5a 1239 993 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.p7b 4535 1239 1400 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b0.p7a 1400 1239 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b0.p10 4535 1242 1105 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b0.p13 1105 1402 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b0.p6c 4535 1240 1241 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b0.p6b 1241 1240 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b0.p6a 4535 1240 1241 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b0.p8c 1241 1402 1242 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b0.p14c 1402 1242 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_b0.p8b 1242 1402 1241 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b0.p18b 4478 1398 1399 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b0.p17c 1398 1278 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.p8a 1241 1402 1242 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b0.p9 1242 4535 1402 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b0.p12 1402 4535 1105 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b0.p5b 4478 993 1239 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.p1 4478 4540 1104 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.p14a 1402 1242 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_b0.p11 1402 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_b0.p18c 1399 1398 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a0.p17d 4478 3572 3660 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.p14d 4535 3453 3662 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_a0.p18f 4478 3660 3661 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a0.p18d 4478 3660 3661 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a0.p2 3406 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.p17a 3660 3572 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.p0 4478 4540 3300 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.p4b 4478 3406 3451 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.p14b 4535 3453 3662 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_a0.p16 3572 3660 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_a0.p17b 4478 3572 3660 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.p4a 3451 3406 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.p18a 3661 3660 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a0.p18e 3661 3660 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a0.p3 3405 3300 3406 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.p7c 3686 3450 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a0.p5a 3450 3405 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.p7b 4535 3450 3686 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a0.p7a 3686 3450 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a0.p10 4535 3453 3452 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a0.p13 3452 3662 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a0.p6c 4535 3451 3454 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a0.p6b 3454 3451 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a0.p6a 4535 3451 3454 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a0.p8c 3454 3662 3453 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a0.p14c 3662 3453 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_a0.p8b 3453 3662 3454 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a0.p18b 4478 3660 3661 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a0.p17c 3660 3572 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.p8a 3454 3662 3453 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a0.p9 3453 4535 3662 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a0.p12 3662 4535 3452 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a0.p5b 4478 3405 3450 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.p1 4478 4540 3406 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.p14a 3662 3453 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_a0.p11 3662 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_a0.p18c 3661 3660 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vsseck1.68onymous_ 4445 4473 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vsseck1.94onymous_ 4473 4476 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vsseck1.25onymous_ 4445 4474 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vsseck1.88onymous_ 4478 4473 4445 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vsseck1.82onymous_ 4445 4473 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vsseck1.77onymous_ 4478 4473 4445 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vsseck1.42onymous_ 4478 4476 4474 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vsseck1.16onymous_ 4478 4474 4445 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vsseck1.36onymous_ 4445 4474 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vsseck1.30onymous_ 4478 4474 4445 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_r3.p18b 4478 4355 4350 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_r3.p17c 4355 4359 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.p1 4478 4368 4367 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.p5b 4478 4373 4374 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.p14a 4371 4370 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_r3.p11 4371 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_r3.p18c 4350 4355 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_r3.p17d 4478 4359 4355 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.p14d 4535 4370 4371 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_r3.p18f 4478 4355 4350 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_r3.p2 4367 4372 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.p18d 4478 4355 4350 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_r3.p17a 4355 4359 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.p4b 4478 4367 4364 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.p0 4478 4372 4375 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.p14b 4535 4370 4371 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_r3.p16 4359 4355 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_r3.p4a 4364 4367 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.p7c 4366 4374 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r3.p17b 4478 4359 4355 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.p7b 4535 4374 4366 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r3.p18a 4350 4355 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_r3.p7a 4366 4374 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r3.p10 4535 4370 4381 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r3.p18e 4350 4355 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_r3.p13 4381 4371 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r3.p3 4373 4375 4367 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.p5a 4374 4373 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.p6c 4535 4364 4365 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r3.p6b 4365 4364 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r3.p6a 4535 4364 4365 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r3.p8c 4365 4371 4370 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r3.p8b 4370 4371 4365 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r3.p8a 4365 4371 4370 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r3.p9 4370 4535 4371 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r3.p12 4371 4535 4381 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r3.p14c 4371 4370 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_q3.p18b 4478 3933 4071 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_q3.p17c 3933 3970 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.p1 4478 4084 4082 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.p5b 4478 4129 4130 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.p14a 4128 4126 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_q3.p11 4128 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_q3.p18c 4071 3933 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_q3.p17d 4478 3970 3933 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.p14d 4535 4126 4128 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_q3.p18f 4478 3933 4071 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_q3.p2 4082 4121 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.p18d 4478 3933 4071 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_q3.p17a 3933 3970 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.p4b 4478 4082 4079 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.p0 4478 4121 4083 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.p14b 4535 4126 4128 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_q3.p16 3970 3933 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_q3.p4a 4079 4082 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.p7c 4081 4130 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q3.p17b 4478 3970 3933 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.p7b 4535 4130 4081 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q3.p18a 4071 3933 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_q3.p7a 4081 4130 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q3.p10 4535 4126 4127 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q3.p18e 4071 3933 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_q3.p13 4127 4128 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q3.p3 4129 4083 4082 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.p5a 4130 4129 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.p6c 4535 4079 4080 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q3.p6b 4080 4079 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q3.p6a 4535 4079 4080 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q3.p8c 4080 4128 4126 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q3.p8b 4126 4128 4080 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q3.p8a 4080 4128 4126 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q3.p9 4126 4535 4128 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q3.p12 4128 4535 4127 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q3.p14c 4128 4126 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_y3.p17d 4478 4417 4418 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.p18c 4419 4418 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y3.p18f 4478 4418 4419 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y3.p14d 4535 4496 4536 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_y3.p18d 4478 4418 4419 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y3.p2 4416 4413 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.p17a 4418 4417 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.p4b 4478 4416 4480 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.p0 4478 4413 4415 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.p16 4417 4418 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_y3.p14b 4535 4496 4536 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_y3.p17b 4478 4417 4418 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.p4a 4480 4416 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.p7c 4498 4479 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y3.p18e 4419 4418 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y3.p7b 4535 4479 4498 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y3.p18a 4419 4418 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y3.p7a 4498 4479 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y3.p10 4535 4496 4495 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y3.p3 4414 4415 4416 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.p13 4495 4536 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y3.p5a 4479 4414 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.p6c 4535 4480 4497 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y3.p6b 4497 4480 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y3.p6a 4535 4480 4497 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y3.p8c 4497 4536 4496 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y3.p8b 4496 4536 4497 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y3.p17c 4418 4417 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.p8a 4497 4536 4496 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y3.p9 4496 4535 4536 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y3.p12 4536 4535 4495 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y3.p14c 4536 4496 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_y3.p18b 4478 4418 4419 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y3.p1 4478 4412 4416 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.p5b 4478 4414 4479 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.p14a 4536 4496 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_y3.p11 4536 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_np.p17a 2754 2860 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.p18d 4478 2754 2717 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_np.p14d 4535 3026 3027 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_np.p18f 4478 2754 2717 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_np.p18c 2717 2754 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_np.p17d 4478 2860 2754 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.p11 3027 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_np.p14a 3027 3026 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_np.p1 4478 3188 2982 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.p12 3027 4535 3137 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_np.p9 3026 4535 3027 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_np.p5b 4478 3028 3030 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.p8a 2980 3027 3026 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_np.p8b 3026 3027 2980 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_np.p8c 2980 3027 3026 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_np.p14c 3027 3026 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_np.p6a 4535 2979 2980 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_np.p18b 4478 2754 2717 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_np.p6b 2980 2979 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_np.p6c 4535 2979 2980 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_np.p17c 2754 2860 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.p13 3137 3027 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_np.p10 4535 3026 3137 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_np.p7a 2981 3030 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_np.p7b 4535 3030 2981 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_np.p7c 2981 3030 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_np.p3 3028 3029 2982 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.p5a 3030 3028 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.p4a 2979 2982 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.p18a 2717 2754 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_np.p18e 2717 2754 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_np.p17b 4478 2860 2754 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.p16 2860 2754 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_np.p14b 4535 3026 3027 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_np.p4b 4478 2982 2979 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.p0 4478 4478 3029 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.p2 2982 4478 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ck.p14a 180 178 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_ck.p18a 4476 172 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_ck.p11 180 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_ck.p17c 172 174 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ck.p18f 4478 172 4476 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_ck.p17a 172 174 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ck.p17d 4478 174 172 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ck.p7c 169 4535 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ck.p18b 4478 172 4476 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_ck.p18e 4476 172 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_ck.p7b 4535 4535 169 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ck.p7a 169 4535 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ck.p10 4535 178 179 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ck.p13 179 180 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ck.p6c 4535 4541 168 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ck.p6b 168 4541 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ck.p14b 4535 178 180 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_ck.p6a 4535 4541 168 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ck.p8c 168 180 178 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ck.p8b 178 180 168 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ck.p8a 168 180 178 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ck.p9 178 4535 180 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ck.p12 180 4535 179 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ck.p16 174 172 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_ck.p18c 4476 172 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_ck.p14c 180 178 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_ck.p18d 4478 172 4476 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_ck.p14d 4535 178 180 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_ck.p17b 4478 174 172 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.p17d 4478 104 105 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.p14d 4535 31 34 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i2.p18f 4478 105 3647 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i2.p18d 4478 105 3647 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i2.p2 101 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.p17a 105 104 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.p0 4478 4540 99 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.p4b 4478 101 102 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.p14b 4535 31 34 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i2.p16 104 105 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_i2.p17b 4478 104 105 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.p4a 102 101 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.p18a 3647 105 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i2.p18e 3647 105 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i2.p3 100 99 101 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.p7c 35 98 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i2.p5a 98 100 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.p7b 4535 98 35 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i2.p7a 35 98 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i2.p10 4535 31 32 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i2.p13 32 34 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i2.p6c 4535 102 33 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i2.p6b 33 102 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i2.p6a 4535 102 33 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i2.p8c 33 34 31 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i2.p14c 34 31 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i2.p8b 31 34 33 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i2.p18b 4478 105 3647 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i2.p17c 105 104 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.p8a 33 34 31 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i2.p9 31 4535 34 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i2.p12 34 4535 32 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i2.p5b 4478 100 98 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.p1 4478 4540 101 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.p14a 34 31 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_i2.p11 34 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_i2.p18c 3647 105 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_f3.p17a 136 139 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.p18d 4478 136 132 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_f3.p14d 4535 150 151 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_f3.p18f 4478 136 132 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_f3.p18c 132 136 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_f3.p17d 4478 139 136 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.p11 151 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_f3.p14a 151 150 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_f3.p1 4478 148 147 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.p12 151 4535 160 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_f3.p9 150 4535 151 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_f3.p5b 4478 152 154 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.p8a 145 151 150 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_f3.p8b 150 151 145 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_f3.p8c 145 151 150 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_f3.p14c 151 150 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_f3.p6a 4535 144 145 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_f3.p18b 4478 136 132 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_f3.p6b 145 144 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_f3.p6c 4535 144 145 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_f3.p17c 136 139 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.p13 160 151 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_f3.p10 4535 150 160 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_f3.p7a 146 154 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_f3.p7b 4535 154 146 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_f3.p7c 146 154 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_f3.p3 152 153 147 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.p5a 154 152 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.p4a 144 147 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.p18a 132 136 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_f3.p18e 132 136 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_f3.p17b 4478 139 136 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.p16 139 136 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_f3.p14b 4535 150 151 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_f3.p4b 4478 147 144 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.p0 4478 4478 153 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.p2 147 4478 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.p17a 996 1106 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.p18d 4478 996 952 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_zero.p14d 4535 1279 1280 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_zero.p18f 4478 996 952 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_zero.p18c 952 996 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_zero.p17d 4478 1106 996 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.p11 1280 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_zero.p14a 1280 1279 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_zero.p1 4478 2790 1246 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.p12 1280 4535 1403 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_zero.p9 1279 4535 1280 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_zero.p5b 4478 1281 1283 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.p8a 1244 1280 1279 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_zero.p8b 1279 1280 1244 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_zero.p8c 1244 1280 1279 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_zero.p14c 1280 1279 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_zero.p6a 4535 1243 1244 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_zero.p18b 4478 996 952 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_zero.p6b 1244 1243 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_zero.p6c 4535 1243 1244 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_zero.p17c 996 1106 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.p13 1403 1280 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_zero.p10 4535 1279 1403 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_zero.p7a 1245 1283 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_zero.p7b 4535 1283 1245 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_zero.p7c 1245 1283 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_zero.p3 1281 1282 1246 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.p5a 1283 1281 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.p4a 1243 1246 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.p18a 952 996 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_zero.p18e 952 996 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_zero.p17b 4478 1106 996 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.p16 1106 996 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_zero.p14b 4535 1279 1280 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_zero.p4b 4478 1246 1243 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.p0 4478 4478 1282 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.p2 1246 4478 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.p17d 4478 96 97 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.p14d 4535 26 29 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i3.p18f 4478 97 130 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i3.p18d 4478 97 130 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i3.p2 93 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.p17a 97 96 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.p0 4478 4540 91 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.p4b 4478 93 92 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.p14b 4535 26 29 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i3.p16 96 97 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_i3.p17b 4478 96 97 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.p4a 92 93 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.p18a 130 97 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i3.p18e 130 97 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i3.p3 94 91 93 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.p7c 30 90 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i3.p5a 90 94 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.p7b 4535 90 30 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i3.p7a 30 90 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i3.p10 4535 26 27 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i3.p13 27 29 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i3.p6c 4535 92 28 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i3.p6b 28 92 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i3.p6a 4535 92 28 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i3.p8c 28 29 26 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i3.p14c 29 26 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i3.p8b 26 29 28 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i3.p18b 4478 97 130 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i3.p17c 97 96 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.p8a 28 29 26 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i3.p9 26 4535 29 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i3.p12 29 4535 27 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i3.p5b 4478 94 90 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.p1 4478 4540 93 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.p14a 29 26 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_i3.p11 29 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_i3.p18c 130 97 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddeck1.55onymous_ 4478 79 126 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddeck1.107nymous_ 126 78 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddeck1.102nymous_ 4478 78 126 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddeck1.41onymous_ 4478 79 126 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddeck1.67onymous_ 4478 4476 79 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddeck1.50onymous_ 126 79 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddeck1.119nymous_ 78 4476 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddeck1.61onymous_ 126 79 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddeck1.93onymous_ 126 78 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddeck1.113nymous_ 4478 78 126 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_r0.p18b 4478 4376 4377 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_r0.p17c 4376 4369 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.p1 4478 4351 4356 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.p5b 4478 4354 4360 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.p14a 4380 4362 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_r0.p11 4380 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_r0.p18c 4377 4376 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_r0.p17d 4478 4369 4376 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.p14d 4535 4362 4380 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_r0.p18f 4478 4376 4377 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_r0.p2 4356 4352 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.p18d 4478 4376 4377 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_r0.p17a 4376 4369 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.p4b 4478 4356 4361 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.p0 4478 4352 4353 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.p14b 4535 4362 4380 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_r0.p16 4369 4376 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_r0.p4a 4361 4356 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.p7c 4378 4360 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r0.p17b 4478 4369 4376 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.p7b 4535 4360 4378 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r0.p18a 4377 4376 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_r0.p7a 4378 4360 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r0.p10 4535 4362 4357 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r0.p18e 4377 4376 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_r0.p13 4357 4380 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r0.p3 4354 4353 4356 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.p5a 4360 4354 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.p6c 4535 4361 4363 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r0.p6b 4363 4361 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r0.p6a 4535 4361 4363 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r0.p8c 4363 4380 4362 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r0.p8b 4362 4380 4363 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r0.p8a 4363 4380 4362 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r0.p9 4362 4535 4380 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r0.p12 4380 4535 4357 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_r0.p14c 4380 4362 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_q0.p18b 4478 4229 4342 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_q0.p17c 4229 4124 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.p1 4478 3931 3968 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.p5b 4478 3932 4076 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.p14a 4125 4077 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_q0.p11 4125 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_q0.p18c 4342 4229 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_q0.p17d 4478 4124 4229 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.p14d 4535 4077 4125 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_q0.p18f 4478 4229 4342 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_q0.p2 3968 4352 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.p18d 4478 4229 4342 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_q0.p17a 4229 4124 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.p4b 4478 3968 4075 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.p0 4478 4352 3930 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.p14b 4535 4077 4125 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_q0.p16 4124 4229 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_q0.p4a 4075 3968 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.p7c 4230 4076 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q0.p17b 4478 4124 4229 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.p7b 4535 4076 4230 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q0.p18a 4342 4229 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_q0.p7a 4230 4076 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q0.p10 4535 4077 3969 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q0.p18e 4342 4229 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_q0.p13 3969 4125 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q0.p3 3932 3930 3968 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.p5a 4076 3932 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.p6c 4535 4075 4078 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q0.p6b 4078 4075 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q0.p6a 4535 4075 4078 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q0.p8c 4078 4125 4077 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q0.p8b 4077 4125 4078 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q0.p8a 4078 4125 4077 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q0.p9 4077 4535 4125 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q0.p12 4125 4535 3969 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_q0.p14c 4125 4077 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_vssick0.34onymous_ 4478 4471 4444 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vssick0.84onymous_ 4444 4472 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vssick0.29onymous_ 4444 4471 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vssick0.79onymous_ 4478 4472 4444 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vssick0.23onymous_ 4478 4471 4444 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vssick0.73onymous_ 4444 4472 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vssick0.43onymous_ 4444 4471 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vssick0.17onymous_ 4471 4476 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vssick0.93onymous_ 4478 4472 4444 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vssick0.67onymous_ 4478 4476 4472 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b3.p17d 4478 149 155 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.p14d 4535 143 159 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_b3.p18f 4478 155 156 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b3.p18d 4478 155 156 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b3.p2 137 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.p17a 155 149 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.p0 4478 4540 134 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.p4b 4478 137 141 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.p14b 4535 143 159 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_b3.p16 149 155 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_b3.p17b 4478 149 155 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.p4a 141 137 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.p18a 156 155 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b3.p18e 156 155 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b3.p3 133 134 137 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.p7c 157 140 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b3.p5a 140 133 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.p7b 4535 140 157 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b3.p7a 157 140 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b3.p10 4535 143 138 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b3.p13 138 159 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b3.p6c 4535 141 142 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b3.p6b 142 141 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b3.p6a 4535 141 142 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b3.p8c 142 159 143 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b3.p14c 159 143 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_b3.p8b 143 159 142 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b3.p18b 4478 155 156 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b3.p17c 155 149 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.p8a 142 159 143 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b3.p9 143 4535 159 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b3.p12 159 4535 138 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b3.p5b 4478 133 140 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.p1 4478 4540 137 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.p14a 159 143 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_b3.p11 159 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_b3.p18c 156 155 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a3.p17d 4478 1826 1940 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.p14d 4535 1691 1941 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_a3.p18f 4478 1940 2930 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a3.p18d 4478 1940 2930 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a3.p2 1661 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.p17a 1940 1826 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.p0 4478 4540 1548 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.p4b 4478 1661 1689 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.p14b 4535 1691 1941 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_a3.p16 1826 1940 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_a3.p17b 4478 1826 1940 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.p4a 1689 1661 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.p18a 2930 1940 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a3.p18e 2930 1940 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a3.p3 1660 1548 1661 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.p7c 1970 1827 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a3.p5a 1827 1660 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.p7b 4535 1827 1970 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a3.p7a 1970 1827 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a3.p10 4535 1691 1690 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a3.p13 1690 1941 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a3.p6c 4535 1689 1692 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a3.p6b 1692 1689 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a3.p6a 4535 1689 1692 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a3.p8c 1692 1941 1691 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a3.p14c 1941 1691 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_a3.p8b 1691 1941 1692 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a3.p18b 4478 1940 2930 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a3.p17c 1940 1826 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.p8a 1692 1941 1691 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a3.p9 1691 4535 1941 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a3.p12 1941 4535 1690 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a3.p5b 4478 1660 1827 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.p1 4478 4540 1661 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.p14a 1941 1691 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_a3.p11 1941 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_a3.p18c 2930 1940 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d2.p17d 4478 4456 4457 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.p14d 4535 4521 4543 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_d2.p18f 4478 4457 4458 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d2.p18d 4478 4457 4458 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d2.p2 4455 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.p17a 4457 4456 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.p0 4478 4540 4453 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.p4b 4478 4455 4489 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.p14b 4535 4521 4543 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_d2.p16 4456 4457 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_d2.p17b 4478 4456 4457 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.p4a 4489 4455 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.p18a 4458 4457 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d2.p18e 4458 4457 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d2.p3 4454 4453 4455 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.p7c 4523 4490 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d2.p5a 4490 4454 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.p7b 4535 4490 4523 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d2.p7a 4523 4490 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d2.p10 4535 4521 4520 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d2.p13 4520 4543 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d2.p6c 4535 4489 4522 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d2.p6b 4522 4489 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d2.p6a 4535 4489 4522 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d2.p8c 4522 4543 4521 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d2.p14c 4543 4521 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_d2.p8b 4521 4543 4522 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d2.p18b 4478 4457 4458 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d2.p17c 4457 4456 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.p8a 4522 4543 4521 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d2.p9 4521 4535 4543 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d2.p12 4543 4535 4520 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d2.p5b 4478 4454 4490 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.p1 4478 4540 4455 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.p14a 4543 4521 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_d2.p11 4543 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_d2.p18c 4458 4457 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i8.p17d 4478 52 53 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.p14d 4535 1 4 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i8.p18f 4478 53 122 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i8.p18d 4478 53 122 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i8.p2 49 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.p17a 53 52 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.p0 4478 4540 48 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.p4b 4478 49 50 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.p14b 4535 1 4 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i8.p16 52 53 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_i8.p17b 4478 52 53 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.p4a 50 49 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.p18a 122 53 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i8.p18e 122 53 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i8.p3 47 48 49 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.p7c 5 46 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i8.p5a 46 47 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.p7b 4535 46 5 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i8.p7a 5 46 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i8.p10 4535 1 2 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i8.p13 2 4 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i8.p6c 4535 50 3 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i8.p6b 3 50 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i8.p6a 4535 50 3 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i8.p8c 3 4 1 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i8.p14c 4 1 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i8.p8b 1 4 3 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i8.p18b 4478 53 122 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i8.p17c 53 52 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.p8a 3 4 1 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i8.p9 1 4535 4 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i8.p12 4 4535 2 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i8.p5b 4478 47 46 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.p1 4478 4540 49 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.p14a 4 1 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_i8.p11 4 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_i8.p18c 122 53 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y1.p17d 4478 4433 4434 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.p18c 4435 4434 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y1.p18f 4478 4434 4435 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y1.p14d 4535 4507 4538 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_y1.p18d 4478 4434 4435 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y1.p2 4432 4430 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.p17a 4434 4433 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.p4b 4478 4432 4483 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.p0 4478 4430 4428 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.p16 4433 4434 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_y1.p14b 4535 4507 4538 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_y1.p17b 4478 4433 4434 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.p4a 4483 4432 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.p7c 4508 4484 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y1.p18e 4435 4434 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y1.p7b 4535 4484 4508 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y1.p18a 4435 4434 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y1.p7a 4508 4484 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y1.p10 4535 4507 4505 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y1.p3 4431 4428 4432 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.p13 4505 4538 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y1.p5a 4484 4431 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.p6c 4535 4483 4506 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y1.p6b 4506 4483 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y1.p6a 4535 4483 4506 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y1.p8c 4506 4538 4507 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y1.p8b 4507 4538 4506 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y1.p17c 4434 4433 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.p8a 4506 4538 4507 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y1.p9 4507 4535 4538 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y1.p12 4538 4535 4505 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y1.p14c 4538 4507 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_y1.p18b 4478 4434 4435 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y1.p1 4478 4429 4432 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.p5b 4478 4431 4484 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.p14a 4538 4507 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_y1.p11 4538 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_vddeck0.55onymous_ 4478 81 127 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddeck0.107nymous_ 127 80 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddeck0.102nymous_ 4478 80 127 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddeck0.41onymous_ 4478 81 127 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddeck0.67onymous_ 4478 4476 81 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddeck0.50onymous_ 127 81 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddeck0.119nymous_ 80 4476 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddeck0.61onymous_ 127 81 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddeck0.93onymous_ 127 80 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddeck0.113nymous_ 4478 80 127 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i4.p17d 4478 88 89 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.p14d 4535 21 24 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i4.p18f 4478 89 128 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i4.p18d 4478 89 128 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i4.p2 85 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.p17a 89 88 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.p0 4478 4540 84 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.p4b 4478 85 86 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.p14b 4535 21 24 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i4.p16 88 89 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_i4.p17b 4478 88 89 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.p4a 86 85 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.p18a 128 89 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i4.p18e 128 89 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i4.p3 83 84 85 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.p7c 25 82 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i4.p5a 82 83 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.p7b 4535 82 25 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i4.p7a 25 82 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i4.p10 4535 21 22 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i4.p13 22 24 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i4.p6c 4535 86 23 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i4.p6b 23 86 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i4.p6a 4535 86 23 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i4.p8c 23 24 21 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i4.p14c 24 21 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i4.p8b 21 24 23 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i4.p18b 4478 89 128 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i4.p17c 89 88 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.p8a 23 24 21 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i4.p9 21 4535 24 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i4.p12 24 4535 22 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i4.p5b 4478 83 82 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.p1 4478 4540 85 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.p14a 24 21 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_i4.p11 24 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_i4.p18c 128 89 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b2.p17d 4478 170 175 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.p14d 4535 166 177 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_b2.p18f 4478 175 176 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b2.p18d 4478 175 176 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b2.p2 163 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.p17a 175 170 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.p0 4478 4540 161 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.p4b 4478 163 164 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.p14b 4535 166 177 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_b2.p16 170 175 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_b2.p17b 4478 170 175 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.p4a 164 163 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.p18a 176 175 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b2.p18e 176 175 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b2.p3 162 161 163 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.p7c 200 171 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b2.p5a 171 162 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.p7b 4535 171 200 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b2.p7a 200 171 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b2.p10 4535 166 165 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b2.p13 165 177 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b2.p6c 4535 164 167 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b2.p6b 167 164 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b2.p6a 4535 164 167 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b2.p8c 167 177 166 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b2.p14c 177 166 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_b2.p8b 166 177 167 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b2.p18b 4478 175 176 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b2.p17c 175 170 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.p8a 167 177 166 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b2.p9 166 4535 177 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b2.p12 177 4535 165 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b2.p5b 4478 162 171 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.p1 4478 4540 163 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.p14a 177 166 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_b2.p11 177 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_b2.p18c 176 175 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_noe.p17d 4478 509 475 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.p14d 4535 736 738 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_noe.p18f 4478 475 431 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_noe.p18d 4478 475 431 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_noe.p2 687 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.p17a 475 509 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.p0 4478 4540 688 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.p4b 4478 687 684 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.p14b 4535 736 738 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_noe.p16 509 475 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_noe.p17b 4478 509 475 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.p4a 684 687 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.p18a 431 475 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_noe.p18e 431 475 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_noe.p3 739 688 687 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.p7c 686 740 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_noe.p5a 740 739 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.p7b 4535 740 686 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_noe.p7a 686 740 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_noe.p10 4535 736 737 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_noe.p13 737 738 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_noe.p6c 4535 684 685 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_noe.p6b 685 684 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_noe.p6a 4535 684 685 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_noe.p8c 685 738 736 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_noe.p14c 738 736 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_noe.p8b 736 738 685 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_noe.p18b 4478 475 431 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_noe.p17c 475 509 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.p8a 685 738 736 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_noe.p9 736 4535 738 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_noe.p12 738 4535 737 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_noe.p5b 4478 739 740 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.p1 4478 4540 687 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.p14a 738 736 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_noe.p11 738 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_noe.p18c 431 475 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_ng.p17a 3407 3408 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.p18d 4478 3407 3235 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_ng.p14d 4535 3663 3573 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_ng.p18f 4478 3407 3235 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_ng.p18c 3235 3407 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_ng.p17d 4478 3408 3407 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.p11 3573 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_ng.p14a 3573 3663 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_ng.p1 4478 3493 3574 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.p12 3573 4535 3664 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ng.p9 3663 4535 3573 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ng.p5b 4478 3576 3575 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.p8a 3455 3573 3663 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ng.p8b 3663 3573 3455 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ng.p8c 3455 3573 3663 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ng.p14c 3573 3663 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_ng.p6a 4535 3457 3455 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ng.p18b 4478 3407 3235 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_ng.p6b 3455 3457 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ng.p6c 4535 3457 3455 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ng.p17c 3407 3408 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.p13 3664 3573 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ng.p10 4535 3663 3664 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ng.p7a 3456 3575 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ng.p7b 4535 3575 3456 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ng.p7c 3456 3575 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_ng.p3 3576 3577 3574 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.p5a 3575 3576 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.p4a 3457 3574 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.p18a 3235 3407 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_ng.p18e 3235 3407 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_ng.p17b 4478 3408 3407 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.p16 3408 3407 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_ng.p14b 4535 3663 3573 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_ng.p4b 4478 3574 3457 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.p0 4478 4478 3577 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.p2 3574 4478 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.p17d 4478 120 121 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.p14d 4535 41 44 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i0.p18f 4478 121 131 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i0.p18d 4478 121 131 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i0.p2 116 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.p17a 121 120 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.p0 4478 4540 115 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.p4b 4478 116 117 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.p14b 4535 41 44 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i0.p16 120 121 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_i0.p17b 4478 120 121 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.p4a 117 116 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.p18a 131 121 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i0.p18e 131 121 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i0.p3 118 115 116 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.p7c 45 114 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i0.p5a 114 118 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.p7b 4535 114 45 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i0.p7a 45 114 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i0.p10 4535 41 42 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i0.p13 42 44 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i0.p6c 4535 117 43 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i0.p6b 43 117 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i0.p6a 4535 117 43 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i0.p8c 43 44 41 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i0.p14c 44 41 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i0.p8b 41 44 43 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i0.p18b 4478 121 131 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i0.p17c 121 120 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.p8a 43 44 41 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i0.p9 41 4535 44 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i0.p12 44 4535 42 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i0.p5b 4478 118 114 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.p1 4478 4540 116 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.p14a 44 41 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_i0.p11 44 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_i0.p18c 131 121 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a1.p17d 4478 3025 3132 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.p14d 4535 2978 3136 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_a1.p18f 4478 3132 3133 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a1.p18d 4478 3132 3133 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a1.p2 2858 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.p17a 3132 3025 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.p0 4478 4540 2752 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.p4b 4478 2858 2976 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.p14b 4535 2978 3136 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_a1.p16 3025 3132 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_a1.p17b 4478 3025 3132 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.p4a 2976 2858 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.p18a 3133 3132 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a1.p18e 3133 3132 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a1.p3 2751 2752 2858 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.p7c 3134 2975 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a1.p5a 2975 2751 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.p7b 4535 2975 3134 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a1.p7a 3134 2975 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a1.p10 4535 2978 2859 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a1.p13 2859 3136 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a1.p6c 4535 2976 2977 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a1.p6b 2977 2976 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a1.p6a 4535 2976 2977 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a1.p8c 2977 3136 2978 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a1.p14c 3136 2978 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_a1.p8b 2978 3136 2977 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a1.p18b 4478 3132 3133 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a1.p17c 3132 3025 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.p8a 2977 3136 2978 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a1.p9 2978 4535 3136 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a1.p12 3136 4535 2859 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a1.p5b 4478 2751 2975 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.p1 4478 4540 2858 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.p14a 3136 2978 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_a1.p11 3136 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_a1.p18c 3133 3132 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b1.p17d 4478 734 819 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.p14d 4535 682 735 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_b1.p18f 4478 819 820 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b1.p18d 4478 819 820 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b1.p2 506 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.p17a 819 734 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.p0 4478 4540 473 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.p4b 4478 506 680 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.p14b 4535 682 735 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_b1.p16 734 819 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_b1.p17b 4478 734 819 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.p4a 680 506 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.p18a 820 819 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b1.p18e 820 819 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b1.p3 474 473 506 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.p7c 821 681 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b1.p5a 681 474 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.p7b 4535 681 821 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b1.p7a 821 681 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b1.p10 4535 682 507 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b1.p13 507 735 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b1.p6c 4535 680 683 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b1.p6b 683 680 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b1.p6a 4535 680 683 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b1.p8c 683 735 682 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b1.p14c 735 682 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_b1.p8b 682 735 683 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b1.p18b 4478 819 820 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_b1.p17c 819 734 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.p8a 683 735 682 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b1.p9 682 4535 735 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b1.p12 735 4535 507 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_b1.p5b 4478 474 681 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.p1 4478 4540 506 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.p14a 735 682 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_b1.p11 735 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_b1.p18c 820 819 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddick0.79onymous_ 4478 2121 2422 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddick0.73onymous_ 2422 2121 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddick0.41onymous_ 2422 2421 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddick0.67onymous_ 4478 4476 2121 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddick0.93onymous_ 4478 2121 2422 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddick0.32onymous_ 4478 2421 2422 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddick0.27onymous_ 2422 2421 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddick0.84onymous_ 2422 2121 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddick0.21onymous_ 4478 2421 2422 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vddick0.15onymous_ 2421 4476 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i5.p17d 4478 76 77 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.p14d 4535 16 19 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i5.p18f 4478 77 125 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i5.p18d 4478 77 125 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i5.p2 73 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.p17a 77 76 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.p0 4478 4540 72 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.p4b 4478 73 74 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.p14b 4535 16 19 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i5.p16 76 77 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_i5.p17b 4478 76 77 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.p4a 74 73 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.p18a 125 77 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i5.p18e 125 77 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i5.p3 71 72 73 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.p7c 20 70 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i5.p5a 70 71 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.p7b 4535 70 20 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i5.p7a 20 70 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i5.p10 4535 16 17 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i5.p13 17 19 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i5.p6c 4535 74 18 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i5.p6b 18 74 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i5.p6a 4535 74 18 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i5.p8c 18 19 16 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i5.p14c 19 16 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i5.p8b 16 19 18 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i5.p18b 4478 77 125 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i5.p17c 77 76 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.p8a 18 19 16 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i5.p9 16 4535 19 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i5.p12 19 4535 17 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i5.p5b 4478 71 70 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.p1 4478 4540 73 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.p14a 19 16 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_i5.p11 19 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_i5.p18c 125 77 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y2.p17d 4478 4425 4426 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.p18c 4427 4426 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y2.p18f 4478 4426 4427 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y2.p14d 4535 4502 4537 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_y2.p18d 4478 4426 4427 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y2.p2 4424 4422 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.p17a 4426 4425 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.p4b 4478 4424 4481 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.p0 4478 4422 4421 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.p16 4425 4426 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_y2.p14b 4535 4502 4537 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_y2.p17b 4478 4425 4426 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.p4a 4481 4424 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.p7c 4503 4482 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y2.p18e 4427 4426 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y2.p7b 4535 4482 4503 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y2.p18a 4427 4426 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y2.p7a 4503 4482 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y2.p10 4535 4502 4500 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y2.p3 4420 4421 4424 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.p13 4500 4537 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y2.p5a 4482 4420 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.p6c 4535 4481 4501 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y2.p6b 4501 4481 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y2.p6a 4535 4481 4501 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y2.p8c 4501 4537 4502 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y2.p8b 4502 4537 4501 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y2.p17c 4426 4425 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.p8a 4501 4537 4502 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y2.p9 4502 4535 4537 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y2.p12 4537 4535 4500 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_y2.p14c 4537 4502 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_y2.p18b 4478 4426 4427 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_y2.p1 4478 4423 4424 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.p5b 4478 4420 4482 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.p14a 4537 4502 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_y2.p11 4537 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_a2.p17d 4478 2466 2573 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.p14d 4535 2419 2467 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_a2.p18f 4478 2573 2929 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a2.p18d 4478 2573 2929 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a2.p2 2282 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.p17a 2573 2466 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.p0 4478 4540 2242 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.p4b 4478 2282 2417 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.p14b 4535 2419 2467 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_a2.p16 2466 2573 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_a2.p17b 4478 2466 2573 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.p4a 2417 2282 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.p18a 2929 2573 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a2.p18e 2929 2573 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a2.p3 2243 2242 2282 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.p7c 2574 2418 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a2.p5a 2418 2243 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.p7b 4535 2418 2574 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a2.p7a 2574 2418 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a2.p10 4535 2419 2283 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a2.p13 2283 2467 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a2.p6c 4535 2417 2420 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a2.p6b 2420 2417 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a2.p6a 4535 2417 2420 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a2.p8c 2420 2467 2419 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a2.p14c 2467 2419 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_a2.p8b 2419 2467 2420 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a2.p18b 4478 2573 2929 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_a2.p17c 2573 2466 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.p8a 2420 2467 2419 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a2.p9 2419 4535 2467 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a2.p12 2467 4535 2283 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_a2.p5b 4478 2243 2418 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.p1 4478 4540 2282 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.p14a 2467 2419 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_a2.p11 2467 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_a2.p18c 2929 2573 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d3.p17d 4478 4450 4451 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.p14d 4535 4516 4542 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_d3.p18f 4478 4451 4452 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d3.p18d 4478 4451 4452 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d3.p2 4449 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.p17a 4451 4450 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.p0 4478 4540 4448 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.p4b 4478 4449 4488 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.p14b 4535 4516 4542 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_d3.p16 4450 4451 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_d3.p17b 4478 4450 4451 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.p4a 4488 4449 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.p18a 4452 4451 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d3.p18e 4452 4451 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d3.p3 4447 4448 4449 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.p7c 4518 4487 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d3.p5a 4487 4447 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.p7b 4535 4487 4518 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d3.p7a 4518 4487 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d3.p10 4535 4516 4515 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d3.p13 4515 4542 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d3.p6c 4535 4488 4517 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d3.p6b 4517 4488 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d3.p6a 4535 4488 4517 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d3.p8c 4517 4542 4516 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d3.p14c 4542 4516 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_d3.p8b 4516 4542 4517 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d3.p18b 4478 4451 4452 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_d3.p17c 4451 4450 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.p8a 4517 4542 4516 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d3.p9 4516 4535 4542 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d3.p12 4542 4535 4515 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_d3.p5b 4478 4447 4487 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.p1 4478 4540 4449 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.p14a 4542 4516 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_d3.p11 4542 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_d3.p18c 4452 4451 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i1.p17d 4478 112 113 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.p14d 4535 36 39 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i1.p18f 4478 113 3559 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i1.p18d 4478 113 3559 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i1.p2 109 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.p17a 113 112 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.p0 4478 4540 108 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.p4b 4478 109 110 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.p14b 4535 36 39 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i1.p16 112 113 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_i1.p17b 4478 112 113 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.p4a 110 109 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.p18a 3559 113 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i1.p18e 3559 113 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i1.p3 107 108 109 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.p7c 40 106 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i1.p5a 106 107 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.p7b 4535 106 40 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i1.p7a 40 106 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i1.p10 4535 36 37 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i1.p13 37 39 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i1.p6c 4535 110 38 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i1.p6b 38 110 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i1.p6a 4535 110 38 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i1.p8c 38 39 36 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i1.p14c 39 36 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i1.p8b 36 39 38 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i1.p18b 4478 113 3559 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i1.p17c 113 112 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.p8a 38 39 36 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i1.p9 36 4535 39 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i1.p12 39 4535 37 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i1.p5b 4478 107 106 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.p1 4478 4540 109 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.p14a 39 36 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_i1.p11 39 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_i1.p18c 3559 113 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vsseck0.68onymous_ 4446 4475 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vsseck0.94onymous_ 4475 4476 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vsseck0.25onymous_ 4446 4477 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vsseck0.88onymous_ 4478 4475 4446 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vsseck0.82onymous_ 4446 4475 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vsseck0.77onymous_ 4478 4475 4446 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vsseck0.42onymous_ 4478 4476 4477 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vsseck0.16onymous_ 4478 4477 4446 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vsseck0.36onymous_ 4446 4477 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_vsseck0.30onymous_ 4478 4477 4446 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_cout.p17a 4388 4389 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.p18d 4478 4388 4382 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_cout.p14d 4535 4399 4400 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_cout.p18f 4478 4388 4382 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_cout.p18c 4382 4388 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_cout.p17d 4478 4389 4388 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.p11 4400 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_cout.p14a 4400 4399 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_cout.p1 4478 4397 4401 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.p12 4400 4535 4409 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cout.p9 4399 4535 4400 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cout.p5b 4478 4403 4402 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.p8a 4394 4400 4399 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cout.p8b 4399 4400 4394 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cout.p8c 4394 4400 4399 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cout.p14c 4400 4399 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_cout.p6a 4535 4396 4394 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cout.p18b 4478 4388 4382 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_cout.p6b 4394 4396 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cout.p6c 4535 4396 4394 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cout.p17c 4388 4389 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.p13 4409 4400 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cout.p10 4535 4399 4409 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cout.p7a 4395 4402 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cout.p7b 4535 4402 4395 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cout.p7c 4395 4402 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cout.p3 4403 4404 4401 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.p5a 4402 4403 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.p4a 4396 4401 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.p18a 4382 4388 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_cout.p18e 4382 4388 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_cout.p17b 4478 4389 4388 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.p16 4389 4388 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_cout.p14b 4535 4399 4400 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_cout.p4b 4478 4401 4396 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.p0 4478 4478 4404 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.p2 4401 4478 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.p17d 4478 68 69 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.p14d 4535 11 14 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i6.p18f 4478 69 124 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i6.p18d 4478 69 124 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i6.p2 65 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.p17a 69 68 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.p0 4478 4540 63 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.p4b 4478 65 66 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.p14b 4535 11 14 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i6.p16 68 69 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_i6.p17b 4478 68 69 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.p4a 66 65 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.p18a 124 69 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i6.p18e 124 69 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i6.p3 64 63 65 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.p7c 15 62 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i6.p5a 62 64 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.p7b 4535 62 15 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i6.p7a 15 62 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i6.p10 4535 11 12 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i6.p13 12 14 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i6.p6c 4535 66 13 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i6.p6b 13 66 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i6.p6a 4535 66 13 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i6.p8c 13 14 11 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i6.p14c 14 11 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_i6.p8b 11 14 13 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i6.p18b 4478 69 124 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_i6.p17c 69 68 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.p8a 13 14 11 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i6.p9 11 4535 14 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i6.p12 14 4535 12 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_i6.p5b 4478 64 62 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.p1 4478 4540 65 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.p14a 14 11 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_i6.p11 14 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_i6.p18c 124 69 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_cin.p17d 4478 4398 4406 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.p14d 4535 4392 4408 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_cin.p18f 4478 4406 4407 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_cin.p18d 4478 4406 4407 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_cin.p2 4386 4540 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.p17a 4406 4398 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.p0 4478 4540 4383 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.p4b 4478 4386 4391 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.p14b 4535 4392 4408 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_cin.p16 4398 4406 4478 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_cin.p17b 4478 4398 4406 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.p4a 4391 4386 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.p18a 4407 4406 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_cin.p18e 4407 4406 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_cin.p3 4385 4383 4386 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.p7c 4410 4390 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cin.p5a 4390 4385 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.p7b 4535 4390 4410 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cin.p7a 4410 4390 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cin.p10 4535 4392 4387 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cin.p13 4387 4408 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cin.p6c 4535 4391 4393 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cin.p6b 4393 4391 4535 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cin.p6a 4535 4391 4393 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cin.p8c 4393 4408 4392 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cin.p14c 4408 4392 4535 4478 tp L=0.32U W=22.6U AS=16.95P AD=16.95P PS=46.7U PD=46.7U 
Mp_cin.p8b 4392 4408 4393 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cin.p18b 4478 4406 4407 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mp_cin.p17c 4406 4398 4478 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.p8a 4393 4408 4392 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cin.p9 4392 4535 4408 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cin.p12 4408 4535 4387 4478 tp L=0.32U W=5.05U AS=3.7875P AD=3.7875P PS=11.6U PD=11.6U 
Mp_cin.p5b 4478 4385 4390 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.p1 4478 4540 4386 4478 tp L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.p14a 4408 4392 4535 4478 tp L=0.32U W=19.15U AS=14.3625P AD=14.3625P PS=39.8U PD=39.8U 
Mp_cin.p11 4408 4541 4535 4478 tp L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mp_cin.p18c 4407 4406 4478 4478 tp L=0.32U W=5.62U AS=4.215P AD=4.215P PS=12.75U PD=12.75U 
Mtr_05276 2595 2593 2594 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05275 2594 2785 2595 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05274 2595 2596 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05273 4540 1564 833 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05272 833 1591 831 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05271 831 830 832 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05270 832 829 1004 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05269 4540 365 211 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05268 4540 1842 1972 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05267 4540 1492 1411 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05266 4540 829 825 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05265 4540 1878 1708 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05264 4540 877 846 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05263 4540 708 381 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05262 4540 2802 2426 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05261 2077 2075 2080 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05260 4540 2196 2078 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05259 2080 2084 2079 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05258 2078 2076 2077 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05257 4540 2079 2092 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05256 744 692 691 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05255 4540 744 745 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05254 691 2782 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05253 1122 1412 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05252 4540 1564 1122 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05251 4540 1975 1122 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05250 1122 1118 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05249 1123 1122 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05248 2590 2783 2591 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05247 4540 2590 2593 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05246 2591 2600 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05245 2111 1488 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05244 4540 1487 2111 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05243 4540 1696 1664 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05242 1664 3905 1697 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05241 1514 1446 1447 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05240 4540 1514 1527 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05239 1447 1516 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05238 1490 1405 1404 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05237 4540 1490 1552 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05236 1404 2284 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05235 302 300 301 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05234 4540 302 328 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05233 301 303 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05232 4540 1705 1668 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05231 1668 2778 1706 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05230 403 401 260 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05229 4540 403 402 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05228 260 404 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05227 1426 1321 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05226 1321 1315 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05225 4540 1318 1321 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05224 4540 1428 2620 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05223 1568 1569 1497 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05222 4540 1568 1710 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05221 1497 1591 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05220 1714 1713 1712 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05219 4540 1714 2004 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05218 1712 1710 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05217 1573 1710 1500 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05216 4540 1573 1730 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05215 1500 1782 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05214 1410 1972 1412 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05213 1412 3226 1410 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05212 1410 1492 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05211 2820 3661 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_05210 2737 2929 2821 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05209 4540 2820 2737 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05208 4540 2929 2931 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05207 2931 3661 2932 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05206 4540 2814 2410 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05205 4540 2825 2414 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05204 4540 2934 1646 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05203 2817 2818 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05202 2818 2929 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05201 4540 3661 2818 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05200 1553 1552 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05199 1553 1551 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05198 4540 1556 1553 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05197 4540 1553 1976 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05196 263 265 262 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05195 4540 263 404 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05194 262 1591 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05193 220 1302 219 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05192 4540 220 238 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05191 219 1564 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05190 583 580 582 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05189 4540 583 605 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05188 582 581 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05187 1566 1565 1494 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05186 4540 1566 1569 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05185 1494 1564 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05184 4540 2447 2542 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05183 2289 2584 2288 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05182 2288 2287 2289 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05181 4540 2285 2288 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05180 2424 2289 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05179 4540 1842 1698 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05178 1698 1834 1699 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05177 1699 1833 1843 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05176 741 694 690 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05175 4540 741 743 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05174 690 689 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05173 206 207 205 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05172 4540 206 510 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05171 205 365 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05170 1116 1110 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05169 4540 1118 1116 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05168 4540 1111 1116 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05167 1116 1835 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05166 4540 803 456 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05165 730 456 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05164 4540 459 730 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05163 4540 211 479 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05162 479 1782 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05161 479 212 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05160 4540 1754 1758 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05159 2635 1758 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05158 4540 1755 2635 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05157 2812 2930 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05156 4540 2817 2812 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05155 2811 2930 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05154 4540 2821 2811 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05153 2924 2930 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05152 4540 2932 2924 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05151 2827 2937 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05150 4540 2821 2827 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05149 4540 2766 2782 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05148 1565 1491 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05147 4540 1407 1491 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05146 1408 1697 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05145 1491 1405 1408 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05144 1493 1413 1414 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05143 4540 1493 1516 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05142 1414 1565 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05141 2137 2139 1994 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05140 4540 2137 2138 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05139 1994 2136 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05138 1294 1296 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05137 1296 1301 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05136 4540 2136 1296 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05135 382 383 228 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05134 4540 382 406 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05133 228 1294 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05132 408 407 268 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05131 4540 408 633 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05130 268 406 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05129 439 438 307 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05128 4540 439 441 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05127 307 633 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05126 1285 1552 1247 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05125 1247 1284 1285 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05124 4540 1288 1247 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05123 1287 1285 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05122 216 213 215 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05121 4540 216 265 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05120 215 1302 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05119 267 264 266 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05118 4540 267 303 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05117 266 265 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05116 4540 2812 2335 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05115 2819 2929 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_05114 2736 3661 2823 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05113 4540 2819 2736 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05112 4540 2809 2337 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05111 235 406 234 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05110 4540 235 385 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05109 234 1591 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05108 1501 1516 1424 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05107 4540 1501 1589 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05106 1424 1591 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05105 423 605 293 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05104 4540 423 658 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05103 293 1782 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05102 1788 1785 1784 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05101 4540 1788 1804 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05100 1784 1782 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05099 4540 1911 2222 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05098 4540 2696 2220 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05097 290 300 289 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05096 4540 290 296 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05095 289 291 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05094 545 1294 546 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05093 4540 545 581 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05092 546 1564 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05091 1974 2778 1973 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05090 4540 1974 2290 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05089 1973 1972 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05088 4540 2781 2695 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05087 4540 2781 2301 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05086 2301 2323 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05085 2301 2620 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05084 2527 2449 2446 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05083 4540 2527 2529 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05082 2446 2445 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05081 899 900 897 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05080 4540 899 898 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05079 897 896 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05078 1920 1919 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05077 4540 2542 1920 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05076 2094 2091 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05075 4540 2220 2094 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05074 1914 1913 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05073 4540 2390 1914 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05072 1923 1922 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05071 4540 2222 1923 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05070 4540 2584 1977 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05069 1977 1837 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05068 1977 1838 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05067 4540 693 524 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05066 524 1412 522 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05065 522 1564 694 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05064 4540 1564 519 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05063 519 693 518 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05062 518 1552 692 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05061 4540 1123 1125 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05060 1125 1150 1124 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05059 1124 1299 1133 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05058 1151 1148 1150 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05057 1150 2171 1151 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05056 1151 1298 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05055 1249 1301 1299 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05054 1299 1298 1249 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05053 1249 1297 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05052 4540 1552 1297 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05051 1297 1564 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05050 1297 1838 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05049 2291 2483 2761 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05048 2761 2476 2291 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05047 2291 2582 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05046 4540 2472 2479 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05045 2479 2471 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05044 2479 2806 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05043 2476 2292 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05042 2292 2290 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05041 4540 2782 2292 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05040 2587 2588 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05039 2588 2806 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05038 4540 2589 2588 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05037 2586 2585 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05036 4540 2584 2586 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05035 2577 2468 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05034 4540 2778 2577 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05033 2724 2783 2785 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05032 2785 3835 2724 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05031 2724 2782 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05030 4540 2598 2599 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05029 2599 2601 2597 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05028 2597 2592 2596 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05027 2602 2620 2601 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05026 2601 2621 2602 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05025 2602 2600 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05024 4540 1591 1419 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05023 1419 1499 1418 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05022 1418 1564 2143 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05021 1000 998 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_05020 998 997 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05019 4540 2620 998 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05018 1009 1032 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_05017 956 1972 1008 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05016 4540 1009 956 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05015 1007 1552 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05014 4540 1004 1007 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05013 4540 2136 1248 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05012 1248 1972 1492 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05011 2781 2779 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05010 4540 2778 2781 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_05009 1290 1411 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05008 1290 1407 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05007 4540 2782 1290 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05006 4540 1290 1288 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05005 4540 1701 1702 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05004 1665 1700 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05003 1666 3905 1665 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05002 1701 1705 1666 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_05001 2286 2782 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_05000 2286 2284 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04999 4540 2290 2286 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04998 4540 2286 2285 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04997 2197 785 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04996 4540 1782 2197 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04995 1707 2138 1847 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04994 1847 1844 1707 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04993 1707 1843 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04992 1625 2217 1528 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04991 1528 2070 1625 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04990 4540 1627 1528 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04989 1624 1625 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04988 436 2217 306 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04987 306 913 436 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04986 4540 440 306 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04985 435 436 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04984 325 2217 324 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04983 324 723 325 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04982 4540 326 324 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04981 320 325 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04980 2218 2217 2095 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04979 2095 2688 2218 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04978 4540 2399 2095 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04977 2215 2218 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04976 4540 543 843 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04975 539 763 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04974 542 541 539 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04973 543 544 542 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04972 4540 227 375 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04971 225 855 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04970 226 224 225 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04969 227 229 226 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04968 4540 2781 2322 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04967 2322 2323 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04966 2322 2325 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04965 918 1096 919 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04964 4540 918 1067 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04963 919 917 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04962 1803 1815 1799 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04961 4540 1803 2087 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04960 1799 1798 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04959 1769 1764 1768 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04958 4540 1769 1798 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04957 1768 1765 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04956 1144 2423 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04955 1144 2513 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04954 4540 1143 1144 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04953 4540 1144 1180 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04952 4540 880 879 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04951 879 877 878 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04950 878 1428 887 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04949 4540 722 629 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04948 629 913 628 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04947 628 2197 888 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04946 4540 1806 1808 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04945 1808 1812 1807 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04944 1807 2696 1809 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04943 4540 1774 1772 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04942 1772 1885 1771 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04941 1771 2357 1789 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04940 4540 1794 1796 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04939 1796 1810 1795 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04938 1795 1911 1797 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04937 4540 1774 1777 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04936 1777 1886 1776 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04935 1776 2656 1790 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04934 2026 2022 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04933 4540 2325 2026 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04932 2011 2423 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04931 2011 2513 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04930 4540 2160 2011 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04929 4540 2011 2041 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04928 4540 2059 2062 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04927 2062 2070 2063 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04926 2063 2197 2064 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04925 4540 1879 1757 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04924 1757 1878 1756 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04923 1756 2437 2035 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04922 4540 2178 2037 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04921 2037 2195 2038 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04920 2038 2447 2179 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04919 4540 1984 1986 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04918 1986 2295 1987 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04917 1987 1985 2130 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04916 1980 1976 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04915 1980 1975 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04914 4540 2290 1980 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04913 4540 1980 1984 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04912 1983 1981 1985 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04911 1985 2516 1983 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04910 1983 1977 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04909 517 515 516 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04908 516 2325 517 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04907 517 521 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04906 2472 1839 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04905 1839 1976 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04904 4540 1835 1839 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04903 4540 2587 2583 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04902 2583 2586 2582 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04901 2582 2581 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04900 4540 2579 2581 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04899 4540 2620 2580 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_04898 2580 2576 4540 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_04897 2579 2577 2578 4541 tn L=0.35U W=2.45U AS=1.8865P AD=1.8865P PS=6.45U PD=6.45U 
Mtr_04896 2578 2806 4540 4541 tn L=0.32U W=2.45U AS=1.8375P AD=1.8375P PS=6.4U PD=6.4U 
Mtr_04895 2580 2806 2579 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_04894 2148 2147 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04893 2148 2143 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04892 4540 2146 2148 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04891 4540 2148 2592 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04890 1013 1002 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04889 4540 1032 953 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04888 953 1000 1002 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04887 954 1007 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04886 4540 1001 955 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04885 1002 1008 954 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04884 955 1116 1002 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04883 4540 1896 1530 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04882 1530 1894 1627 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04881 4540 441 313 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04880 313 763 440 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04879 4540 328 327 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04878 327 855 326 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04877 4540 2699 2398 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04876 2398 2457 2399 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04875 4540 1895 1773 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04874 1773 1894 2191 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04873 4540 846 847 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04872 847 2297 845 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04871 845 843 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04870 4540 381 223 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04869 223 2297 380 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04868 380 375 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04867 4540 2426 2298 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04866 2298 2297 2774 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04865 2774 2301 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04864 4540 1885 1747 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04863 4540 1051 696 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04862 4540 2320 2319 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04861 2319 2315 2317 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04860 2317 2322 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04859 1197 1235 1194 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04858 4540 1197 1193 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04857 1194 1192 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04856 1178 1175 1177 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04855 4540 1178 1192 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04854 1177 1176 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04853 873 871 872 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04852 4540 873 917 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04851 872 874 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04850 4540 1072 978 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04849 978 1090 979 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04848 979 1911 1066 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04847 4540 903 902 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04846 902 904 901 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04845 901 2447 900 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04844 4540 714 570 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04843 570 1160 571 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04842 571 2435 896 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04841 4540 1072 975 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04840 975 1061 974 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04839 974 2656 1062 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04838 4540 1809 1793 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04837 1793 1789 1792 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04836 1792 1797 1791 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04835 1791 1790 2202 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04834 4540 2044 2049 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04833 2049 2041 2047 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04832 2047 2042 2048 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04831 2048 2043 2203 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04830 2031 2032 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04829 4540 2513 2031 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04828 2294 2307 2295 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04827 2295 2325 2294 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04826 2294 2516 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04825 4540 2055 2008 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04824 4540 614 604 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04823 604 763 603 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04822 4540 296 287 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04821 287 855 288 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04820 4540 2699 2369 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04819 2369 2544 2366 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04818 4540 1472 1473 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04817 1473 1894 1642 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04816 4540 1347 859 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04815 4540 2356 2320 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04814 4540 1849 1846 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04813 1894 1846 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04812 4540 1847 1894 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04811 761 698 697 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04810 4540 761 763 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04809 697 1287 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04808 1302 1303 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04807 1303 1301 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04806 4540 2284 1303 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04805 4540 1706 1703 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04804 1703 2782 1704 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04803 1704 1702 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04802 849 848 850 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04801 4540 849 855 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04800 850 1704 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04799 2617 2513 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04798 4540 2781 2617 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04797 4540 1851 1711 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04796 1711 1999 2297 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04795 549 581 548 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04794 4540 549 544 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04793 548 1591 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04792 222 238 221 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04791 4540 222 229 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04790 221 1591 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04789 4540 2656 2171 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04788 1590 1589 1511 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04787 4540 1590 1750 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04786 1511 1782 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04785 384 763 232 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04784 4540 384 537 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04783 232 1782 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04782 405 404 261 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04781 4540 405 576 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04780 261 1782 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04779 2657 2695 2658 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04778 4540 2657 2655 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04777 2658 2656 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04776 4540 2357 2325 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04775 4540 1415 1416 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04774 1416 1421 2315 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04773 231 229 230 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04772 4540 231 856 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04771 230 1782 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04770 1111 1108 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04769 1108 1126 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04768 4540 2782 1108 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04767 4540 2034 1882 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04766 4540 2924 2175 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04765 4540 1893 2229 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04764 209 1591 208 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04763 4540 209 693 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04762 208 207 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04761 207 210 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04760 4540 212 207 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04759 4540 1044 521 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04758 827 825 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04757 827 828 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04756 4540 826 827 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04755 4540 827 1838 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04754 1975 1115 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04753 1115 1117 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04752 4540 1111 1115 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04751 4540 2589 2783 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04750 4540 2488 2600 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04749 386 401 233 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04748 4540 386 555 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04747 233 385 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04746 1503 1499 1425 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04745 4540 1503 1862 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04744 1425 1589 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04743 4540 2435 2513 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04742 1040 1024 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04741 1024 1026 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04740 4540 1564 1024 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04739 2481 2424 2425 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04738 4540 2481 2841 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04737 2425 2423 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04736 852 1704 851 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04735 4540 852 853 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04734 851 2423 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04733 764 1287 699 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04732 4540 764 765 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04731 699 2423 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04730 2002 1709 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04729 4540 1847 2002 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04728 2693 2695 2692 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04727 4540 2693 2694 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04726 2692 2691 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04725 294 291 292 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04724 4540 294 332 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04723 292 1782 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04722 2698 2695 2697 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04721 4540 2698 2840 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04720 2697 2696 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04719 304 303 305 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04718 4540 304 661 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04717 305 1782 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04716 635 633 634 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04715 4540 635 728 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04714 634 1782 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04713 1529 1527 1464 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04712 4540 1529 1472 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04711 1464 1782 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04710 2544 2542 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04709 4540 2781 2544 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04708 241 264 240 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04707 4540 241 291 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04706 240 238 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04705 612 608 611 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04704 4540 612 614 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04703 611 605 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04702 1780 1778 1779 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04701 4540 1780 1895 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04700 1779 1785 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04699 1570 1572 1498 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04698 4540 1570 1785 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04697 1498 1569 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04696 1598 1593 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04695 1593 1592 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04694 4540 1591 1593 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04693 4540 2323 2699 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04692 4540 2122 2123 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04691 2584 2123 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04690 4540 4350 2584 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04689 2457 2390 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04688 4540 2781 2457 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04687 2447 1598 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04686 4540 1782 2447 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04685 1521 1458 1456 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04684 4540 1521 2360 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04683 1456 1522 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04682 2696 783 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04681 4540 785 2696 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04680 2120 2117 2119 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04679 4540 2120 2702 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04678 2119 2118 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04677 1911 1460 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04676 4540 1598 1911 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04675 805 731 732 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04674 4540 805 2227 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04673 732 803 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04672 4540 1532 1470 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04671 2455 1470 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04670 4540 1468 2455 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04669 4540 1522 1457 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04668 2199 1457 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04667 4540 1458 2199 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04666 4540 2118 2114 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04665 2844 2114 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04664 4540 2117 2844 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04663 2435 1040 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04662 4540 1782 2435 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04661 2016 2022 2017 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04660 4540 2016 2429 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04659 2017 2020 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04658 1428 1426 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04657 4540 1782 1428 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04656 2656 1038 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04655 4540 1040 2656 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04654 1596 1595 1515 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04653 4540 1596 2352 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04652 1515 1754 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04651 2357 1319 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04650 4540 1426 2357 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04649 4540 2020 2021 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04648 2613 2021 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04647 4540 2022 2613 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04646 4540 363 365 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04645 365 367 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04644 365 1972 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04643 4540 1421 1423 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04642 1585 1423 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04641 4540 1420 1585 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04640 2809 2930 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04639 4540 2823 2809 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04638 2814 2937 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04637 4540 2817 2814 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04636 2825 2937 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04635 4540 2823 2825 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04634 2934 2937 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04633 4540 2932 2934 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04632 4540 2307 2296 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04631 2296 2424 2323 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04630 829 824 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04629 4540 823 829 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04628 1999 2111 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04627 4540 2620 1999 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04626 1421 2111 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04625 4540 2325 1421 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04624 1754 2111 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04623 4540 2171 1754 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04622 2020 2111 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04621 4540 2513 2020 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04620 803 988 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04619 4540 2222 803 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04618 2118 2111 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04617 4540 2220 2118 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04616 1522 2111 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04615 4540 2542 1522 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04614 1532 2111 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04613 4540 2390 1532 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04612 4540 367 1564 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04611 4540 1571 1835 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04610 4540 1126 2423 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04609 4540 520 1591 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04608 4540 3226 1407 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04607 4540 3905 2136 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04606 4540 3911 2284 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04605 4540 3835 2778 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04604 4540 2930 2937 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04603 4540 703 705 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04602 705 704 785 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04601 4540 2197 2390 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04600 1526 1462 1463 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04599 4540 1526 1896 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04598 1463 1527 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04597 1531 1465 1466 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04596 4540 1531 2217 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04595 1466 1532 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04594 1523 1623 1617 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04593 4540 2070 1523 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04592 1617 1621 1615 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04591 4540 1615 1524 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04590 1524 1621 1620 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04589 1620 1623 1525 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04588 1621 1623 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04587 4540 1622 1623 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04586 1525 1618 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04585 4540 1624 1618 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04584 2070 1617 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04583 4540 1617 2070 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04582 1615 1620 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04581 295 433 424 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04580 4540 913 295 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04579 424 434 426 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04578 4540 426 298 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04577 298 434 428 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04576 428 433 299 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04575 434 433 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04574 4540 432 433 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04573 299 429 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04572 4540 435 429 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04571 913 424 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04570 4540 424 913 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04569 426 428 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04568 308 321 310 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04567 4540 723 308 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04566 310 317 309 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04565 4540 309 311 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04564 311 317 312 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04563 312 321 318 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04562 317 321 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04561 4540 314 321 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04560 318 315 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04559 4540 320 315 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04558 723 310 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04557 4540 310 723 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04556 309 312 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04555 2086 2216 2208 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04554 4540 2688 2086 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04553 2208 2210 2209 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04552 4540 2209 2085 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04551 2085 2210 2213 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04550 2213 2216 2090 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04549 2210 2216 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04548 4540 2214 2216 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04547 2090 2211 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04546 4540 2215 2211 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04545 2688 2208 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04544 4540 2208 2688 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04543 2209 2213 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04542 2192 2360 2058 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04541 2058 2195 2192 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04540 4540 2191 2058 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04539 2189 2192 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04538 2045 2190 2183 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04537 4540 2195 2045 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04536 2183 2184 2180 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04535 4540 2180 2046 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04534 2046 2184 2187 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04533 2187 2190 2053 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04532 2184 2190 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04531 4540 2188 2190 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04530 2053 2185 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04529 4540 2189 2185 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04528 2195 2183 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04527 4540 2183 2195 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04526 2180 2187 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04525 601 2360 602 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04524 602 904 601 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04523 4540 603 602 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04522 600 601 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04521 586 599 589 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04520 4540 904 586 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04519 589 598 593 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04518 4540 593 590 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04517 590 598 591 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04516 591 599 592 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04515 598 599 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04514 4540 594 599 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04513 592 597 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04512 4540 600 597 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04511 904 589 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04510 4540 589 904 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04509 593 591 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04508 284 2360 285 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04507 285 715 284 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04506 4540 288 285 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04505 283 284 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04504 270 278 271 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04503 4540 715 270 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04502 271 280 272 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04501 4540 272 276 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04500 276 280 275 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04499 275 278 273 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04498 280 278 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04497 4540 277 278 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04496 273 274 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04495 4540 283 274 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04494 715 271 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04493 4540 271 715 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04492 272 275 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04491 2363 2360 2365 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04490 2365 2826 2363 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04489 4540 2366 2365 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04488 2538 2363 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04487 2364 2533 2535 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04486 4540 2826 2364 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04485 2535 2532 2537 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04484 4540 2537 2367 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04483 2367 2532 2534 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04482 2534 2533 2368 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04481 2532 2533 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04480 4540 2451 2533 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04479 2368 2541 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04478 4540 2538 2541 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04477 2826 2535 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04476 4540 2535 2826 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04475 2537 2534 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04474 1643 2702 1540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04473 1540 1812 1643 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04472 4540 1642 1540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04471 1651 1643 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04470 1544 1658 1650 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04469 4540 1812 1544 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04468 1650 1659 1652 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04467 4540 1652 1546 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04466 1546 1659 1654 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04465 1654 1658 1545 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04464 1659 1658 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04463 4540 1656 1658 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04462 1545 1657 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04461 4540 1651 1657 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04460 1812 1650 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04459 4540 1650 1812 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04458 1652 1654 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04457 4540 728 727 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04456 727 763 1084 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04455 1085 2702 987 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04454 987 1091 1085 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04453 4540 1084 987 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04452 1082 1085 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04451 984 1083 1074 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04450 4540 1091 984 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04449 1074 1080 1075 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04448 4540 1075 985 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04447 985 1080 1078 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04446 1078 1083 986 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04445 1080 1083 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04444 4540 1081 1083 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04443 986 1077 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04442 4540 1082 1077 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04441 1091 1074 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04440 4540 1074 1091 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04439 1075 1078 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04438 4540 661 660 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04437 660 855 1379 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04436 1380 2702 1274 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04435 1274 1382 1380 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04434 4540 1379 1274 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04433 1385 1380 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04432 1275 1394 1384 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04431 4540 1382 1275 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04430 1384 1393 1386 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04429 4540 1386 1276 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04428 1276 1393 1389 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04427 1389 1394 1277 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04426 1393 1394 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04425 4540 1391 1394 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04424 1277 1392 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04423 4540 1385 1392 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04422 1382 1384 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04421 4540 1384 1382 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04420 1386 1389 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04419 4540 2699 2700 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04418 2700 2840 2701 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04417 2704 2702 2703 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04416 2703 2705 2704 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04415 4540 2701 2703 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04414 2708 2704 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04413 2707 2716 2706 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04412 4540 2705 2707 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04411 2706 2715 2709 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04410 4540 2709 2711 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04409 2711 2715 2710 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04408 2710 2716 2712 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04407 2715 2716 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04406 4540 2713 2716 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04405 2712 2714 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04404 4540 2708 2714 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04403 2705 2706 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04402 4540 2706 2705 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04401 2709 2710 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04400 4540 1804 1538 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04399 1538 1894 1641 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04398 1639 2227 1537 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04397 1537 1810 1639 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04396 4540 1641 1537 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04395 1638 1639 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04394 1533 1637 1630 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04393 4540 1810 1533 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04392 1630 1631 1628 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04391 4540 1628 1534 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04390 1534 1631 1635 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04389 1635 1637 1535 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04388 1631 1637 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04387 4540 1636 1637 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04386 1535 1632 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04385 4540 1638 1632 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04384 1810 1630 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04383 4540 1630 1810 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04382 1628 1635 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04381 4540 658 329 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04380 329 763 452 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04379 453 2227 333 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04378 333 1090 453 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04377 4540 452 333 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04376 455 453 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04375 319 449 444 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04374 4540 1090 319 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04373 444 451 445 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04372 4540 445 322 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04371 322 451 447 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04370 447 449 323 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04369 451 449 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04368 4540 448 449 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04367 323 450 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04366 4540 455 450 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04365 1090 444 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04364 4540 444 1090 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04363 445 447 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04362 4540 332 331 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04361 331 855 335 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04360 336 2227 338 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04359 338 1371 336 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04358 4540 335 338 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04357 342 336 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04356 340 351 341 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04355 4540 1371 340 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04354 341 350 343 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04353 4540 343 346 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04352 346 350 348 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04351 348 351 347 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04350 350 351 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04349 4540 349 351 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04348 347 352 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04347 4540 342 352 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04346 1371 341 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04345 4540 341 1371 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04344 343 348 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04343 4540 2699 2400 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04342 2400 2694 2401 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04341 2225 2227 2109 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04340 2109 2677 2225 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04339 4540 2401 2109 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04338 2233 2225 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04337 2113 2240 2232 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04336 4540 2677 2113 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04335 2232 2241 2234 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04334 4540 2234 2115 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04333 2115 2241 2237 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04332 2237 2240 2116 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04331 2241 2240 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04330 4540 2238 2240 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04329 2116 2239 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04328 4540 2233 2239 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04327 2677 2232 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04326 4540 2232 2677 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04325 2234 2237 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04324 4540 1896 1775 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04323 1775 2002 2096 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04322 2097 2099 2098 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04321 2098 2455 2097 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04320 4540 2096 2098 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04319 2106 2097 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04318 2100 2112 2104 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04317 4540 2099 2100 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04316 2104 2108 2101 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04315 4540 2101 2102 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04314 2102 2108 2103 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04313 2103 2112 2110 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04312 2108 2112 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04311 4540 2105 2112 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04310 2110 2107 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04309 4540 2106 2107 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04308 2099 2104 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04307 4540 2104 2099 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04306 2101 2103 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04305 4540 441 316 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04304 316 765 649 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04303 653 926 655 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04302 655 2455 653 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04301 4540 649 655 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04300 651 653 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04299 636 647 637 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04298 4540 926 636 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04297 637 646 640 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04296 4540 640 642 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04295 642 646 641 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04294 641 647 643 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04293 646 647 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04292 4540 644 647 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04291 643 648 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04290 4540 651 648 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04289 926 637 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04288 4540 637 926 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04287 640 641 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04286 4540 328 330 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04285 330 853 654 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04284 657 1206 656 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04283 656 2455 657 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04282 4540 654 656 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04281 796 657 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04280 645 788 791 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04279 4540 1206 645 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04278 791 787 794 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04277 4540 794 652 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04276 652 787 792 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04275 792 788 650 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04274 787 788 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04273 4540 726 788 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04272 650 799 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04271 4540 796 799 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04270 1206 791 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04269 4540 791 1206 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04268 794 792 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04267 4540 2457 2458 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04266 2458 2841 2459 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04265 2555 2684 2393 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04264 2393 2455 2555 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04263 4540 2459 2393 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04262 2556 2555 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04261 2381 2548 2552 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04260 4540 2684 2381 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04259 2552 2546 2551 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04258 4540 2551 2383 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04257 2383 2546 2549 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04256 2549 2548 2387 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04255 2546 2548 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04254 4540 2454 2548 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04253 2387 2554 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04252 4540 2556 2554 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04251 2684 2552 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04250 4540 2552 2684 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04249 2551 2549 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04248 4540 1895 1681 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04247 1681 2002 1897 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04246 1899 2065 1781 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04245 1781 2199 1899 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04244 4540 1897 1781 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04243 1906 1899 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04242 1783 1909 1902 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04241 4540 2065 1783 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04240 1902 1910 1903 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04239 4540 1903 1787 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04238 1787 1910 1905 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04237 1905 1909 1786 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04236 1910 1909 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04235 4540 1907 1909 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04234 1786 1908 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04233 4540 1906 1908 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04232 2065 1902 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04231 4540 1902 2065 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04230 1903 1905 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04229 4540 614 613 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04228 613 765 630 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04227 632 1063 631 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04226 631 2199 632 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04225 4540 630 631 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04224 626 632 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04223 615 627 617 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04222 4540 1063 615 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04221 617 624 616 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04220 4540 616 621 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04219 621 624 622 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04218 622 627 623 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04217 624 627 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04216 4540 625 627 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04215 623 620 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04214 4540 626 620 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04213 1063 617 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04212 4540 617 1063 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04211 616 622 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04210 4540 296 297 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04209 297 853 1200 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04208 1201 1357 1202 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04207 1202 2199 1201 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04206 4540 1200 1202 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04205 1363 1201 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04204 1267 1367 1361 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04203 4540 1357 1267 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04202 1361 1366 1358 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04201 4540 1358 1268 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04200 1268 1366 1360 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04199 1360 1367 1269 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04198 1366 1367 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04197 4540 1362 1367 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04196 1269 1364 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04195 4540 1363 1364 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04194 1357 1361 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04193 4540 1361 1357 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04192 1358 1360 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04191 4540 2544 2452 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04190 2452 2841 2453 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04189 2200 2664 2074 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04188 2074 2199 2200 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04187 4540 2453 2074 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04186 2372 2200 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04185 2371 2380 2370 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04184 4540 2664 2371 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04183 2370 2379 2373 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04182 4540 2373 2375 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04181 2375 2379 2377 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04180 2377 2380 2376 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04179 2379 2380 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04178 4540 2378 2380 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04177 2376 2374 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04176 4540 2372 2374 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04175 2664 2370 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04174 4540 2370 2664 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04173 2373 2377 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04172 4540 1472 1471 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04171 1471 2002 1474 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04170 1539 1915 1476 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04169 1476 2844 1539 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04168 4540 1474 1476 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04167 1478 1539 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04166 1477 1486 1541 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04165 4540 1915 1477 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04164 1541 1485 1543 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04163 4540 1543 1481 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04162 1481 1485 1542 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04161 1542 1486 1482 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04160 1485 1486 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04159 4540 1484 1486 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04158 1482 1483 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04157 4540 1478 1483 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04156 1915 1541 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04155 4540 1541 1915 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04154 1543 1542 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04153 4540 728 729 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04152 729 765 934 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04151 935 1092 936 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04150 936 2844 935 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04149 4540 934 936 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04148 943 935 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04147 942 951 941 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04146 4540 1092 942 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04145 941 950 944 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04144 4540 944 946 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04143 946 950 945 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04142 945 951 947 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04141 950 951 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04140 4540 948 951 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04139 947 949 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04138 4540 943 949 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04137 1092 941 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04136 4540 941 1092 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04135 944 945 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04134 4540 661 663 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04133 663 853 937 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04132 940 1226 939 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04131 939 2844 940 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04130 4540 937 939 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04129 938 940 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04128 668 808 809 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04127 4540 1226 668 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04126 809 807 812 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04125 4540 812 674 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04124 674 807 813 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04123 813 808 675 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04122 807 808 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04121 4540 733 808 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04120 675 818 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04119 4540 938 818 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04118 1226 809 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04117 4540 809 1226 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04116 812 813 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04115 4540 2840 2746 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04114 2746 2841 2842 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04113 2843 2846 2747 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04112 2747 2844 2843 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04111 4540 2842 2747 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04110 2850 2843 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04109 2748 2857 2848 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04108 4540 2846 2748 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04107 2848 2856 2849 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04106 4540 2849 2749 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04105 2749 2856 2853 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04104 2853 2857 2750 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04103 2856 2857 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04102 4540 2854 2857 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04101 2750 2855 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04100 4540 2850 2855 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04099 2846 2848 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04098 4540 2848 2846 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04097 2849 2853 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04096 4540 1804 1682 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04095 1682 2002 1925 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04094 1926 1928 1818 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04093 1818 2463 1926 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04092 4540 1925 1818 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04091 1931 1926 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04090 1820 1937 1930 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04089 4540 1928 1820 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04088 1930 1938 1932 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04087 4540 1932 1822 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04086 1822 1938 1935 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04085 1935 1937 1823 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04084 1938 1937 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04083 4540 1936 1937 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04082 1823 1939 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04081 4540 1931 1939 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04080 1928 1930 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04079 4540 1930 1928 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04078 1932 1935 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04077 4540 658 659 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04076 659 765 662 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04075 665 1095 664 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04074 664 730 665 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04073 4540 662 664 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04072 669 665 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04071 666 678 667 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04070 4540 1095 666 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04069 667 677 670 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04068 4540 670 671 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04067 671 677 673 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04066 673 678 672 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04065 677 678 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04064 4540 676 678 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04063 672 679 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04062 4540 669 679 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04061 1095 667 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04060 4540 667 1095 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04059 670 673 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04058 4540 332 334 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04057 334 853 458 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04056 461 1232 337 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04055 337 730 461 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04054 4540 458 337 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04053 464 461 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04052 339 471 463 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04051 4540 1232 339 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04050 463 472 465 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04049 4540 465 344 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04048 344 472 468 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04047 468 471 345 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04046 472 471 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04045 4540 469 471 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04044 345 470 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04043 4540 464 470 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04042 1232 463 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04041 4540 463 1232 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04040 465 468 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04039 4540 2694 2461 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04038 2461 2841 2462 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04037 2557 2561 2407 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04036 2407 2463 2557 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04035 4540 2462 2407 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04034 2566 2557 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04033 2409 2560 2562 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04032 4540 2561 2409 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04031 2562 2559 2565 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04030 4540 2565 2412 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04029 2412 2559 2567 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04028 2567 2560 2413 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04027 2559 2560 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04026 4540 2465 2560 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04025 2413 2572 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04024 4540 2566 2572 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04023 2561 2562 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04022 4540 2562 2561 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04021 2565 2567 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_04020 1512 1441 1444 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04019 1444 2635 1512 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04018 4540 1438 1444 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04017 1440 1512 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_04016 4540 576 579 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04015 579 853 1438 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04014 1127 1137 1128 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04013 4540 1298 1127 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04012 1128 1136 1129 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04011 4540 1129 1131 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04010 1131 1136 1130 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04009 1130 1137 1132 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04008 1136 1137 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04007 4540 1134 1137 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04006 1132 1135 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04005 4540 1133 1135 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_04004 1298 1128 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04003 4540 1128 1298 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_04002 1129 1130 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_04001 1746 1876 1869 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_04000 4540 2023 1746 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03999 1869 1877 1868 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03998 4540 1868 1748 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03997 1748 1877 1874 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03996 1874 1876 1749 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03995 1877 1876 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03994 4540 1875 1876 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03993 1749 1872 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03992 4540 1870 1872 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03991 2023 1869 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03990 4540 1869 2023 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03989 1868 1874 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03988 1752 2023 1753 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03987 1753 2635 1752 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03986 4540 1751 1753 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03985 1870 1752 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03984 4540 1750 1677 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03983 1677 2002 1751 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03982 2718 2762 2756 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03981 4540 2806 2718 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03980 2756 2765 2757 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03979 4540 2757 2719 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03978 2719 2765 2759 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03977 2759 2762 2720 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03976 2765 2762 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03975 4540 2760 2762 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03974 2720 2763 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03973 4540 2761 2763 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03972 2806 2756 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03971 4540 2756 2806 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03970 2757 2759 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03969 4540 2806 2293 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03968 2293 3911 2483 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03967 2483 2479 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03966 2299 2486 2490 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03965 4540 2488 2299 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03964 2490 2485 2491 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03963 4540 2491 2302 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_03962 2302 2485 2487 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03961 2487 2486 2300 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03960 2485 2486 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03959 4540 2427 2486 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03958 2300 2494 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03957 4540 2594 2494 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03956 2488 2490 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03955 4540 2490 2488 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03954 2491 2487 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_03953 2141 2139 2000 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03952 2000 3911 2141 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03951 4540 2140 2000 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03950 2147 2141 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03949 4540 2138 2140 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03948 957 1021 1012 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03947 4540 1032 957 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03946 1012 1014 1011 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03945 4540 1011 959 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03944 959 1014 1016 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03943 1016 1021 958 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03942 1014 1021 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03941 4540 1020 1021 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03940 958 1015 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03939 4540 1013 1015 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03938 1032 1012 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03937 4540 1012 1032 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03936 1011 1016 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03935 4540 1412 1001 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03934 1989 1997 1988 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03933 4540 2055 1989 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03932 1988 1996 1990 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03931 4540 1990 1991 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03930 1991 1996 1993 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03929 1993 1997 1992 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03928 1996 1997 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03927 4540 1995 1997 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03926 1992 1998 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03925 4540 2005 1998 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03924 2055 1988 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03923 4540 1988 2055 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03922 1990 1993 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03921 2006 2001 4540 4541 tn L=0.35U W=2.45U AS=1.8865P AD=1.8865P PS=6.45U PD=6.45U 
Mtr_03920 2007 2002 4540 4541 tn L=0.32U W=2.45U AS=1.8375P AD=1.8375P PS=6.4U PD=6.4U 
Mtr_03919 4540 2003 2006 4541 tn L=0.35U W=2.45U AS=1.8865P AD=1.8865P PS=6.45U PD=6.45U 
Mtr_03918 2006 2008 2005 4541 tn L=0.35U W=2.45U AS=1.8865P AD=1.8865P PS=6.45U PD=6.45U 
Mtr_03917 2005 2004 2007 4541 tn L=0.35U W=2.45U AS=1.8865P AD=1.8865P PS=6.45U PD=6.45U 
Mtr_03916 4540 1999 2003 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03915 2603 2611 2604 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03914 4540 2801 2603 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03913 2604 2610 2605 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03912 4540 2605 2608 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03911 2608 2610 2607 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03910 2607 2611 2606 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03909 2610 2611 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03908 4540 2609 2611 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03907 2606 2612 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03906 4540 2614 2612 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03905 2801 2604 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03904 4540 2604 2801 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03903 2605 2607 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03902 2615 2801 2616 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03901 2616 2613 2615 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03900 4540 2619 2616 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03899 2614 2615 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03898 4540 2617 2618 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03897 2618 2841 2619 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03896 559 567 564 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03895 4540 1326 559 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03894 564 569 563 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03893 4540 563 565 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03892 565 569 561 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03891 561 567 562 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03890 569 567 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03889 4540 566 567 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03888 562 568 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03887 4540 573 568 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03886 1326 564 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03885 4540 564 1326 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03884 563 561 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03883 4540 1862 1729 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03882 1729 1894 2012 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03881 2015 2429 2014 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03880 2014 2161 2015 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03879 4540 2012 2014 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03878 2153 2015 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03877 2009 2159 2151 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03876 4540 2161 2009 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03875 2151 2154 2149 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03874 4540 2149 2010 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_03873 2010 2154 2157 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03872 2157 2159 2013 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03871 2154 2159 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03870 4540 2158 2159 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03869 2013 2155 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03868 4540 2153 2155 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03867 2161 2151 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03866 4540 2151 2161 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03865 2149 2157 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_03864 4540 555 552 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03863 552 763 553 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03862 550 2429 554 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03861 554 1160 550 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03860 4540 553 554 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03859 547 550 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03858 523 536 529 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03857 4540 1160 523 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03856 529 535 528 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03855 4540 528 530 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_03854 530 535 527 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03853 527 536 526 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03852 535 536 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03851 4540 531 536 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03850 526 533 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03849 4540 547 533 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03848 1160 529 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03847 4540 529 1160 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03846 528 527 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_03845 4540 402 254 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03844 254 855 400 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03843 398 2429 252 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03842 252 1152 398 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03841 4540 400 252 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03840 397 398 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03839 237 396 388 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03838 4540 1152 237 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03837 388 395 389 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03836 4540 389 239 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03835 239 395 391 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03834 391 396 243 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03833 395 396 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03832 4540 392 396 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03831 243 393 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03830 4540 397 393 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03829 1152 388 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03828 4540 388 1152 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03827 389 391 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03826 4540 2699 2431 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03825 2431 2617 2432 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03824 2510 2429 2321 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03823 2321 2497 2510 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03822 4540 2432 2321 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03821 2511 2510 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03820 2314 2499 2502 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03819 4540 2497 2314 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03818 2502 2498 2503 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03817 4540 2503 2318 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03816 2318 2498 2500 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03815 2500 2499 2316 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03814 2498 2499 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03813 4540 2428 2499 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03812 2316 2507 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03811 4540 2511 2507 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03810 2497 2502 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03809 4540 2502 2497 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03808 2503 2500 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03807 1495 1894 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03806 1718 2004 1495 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03805 1496 1708 1718 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03804 4540 2297 1496 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03803 1717 1728 1716 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03802 4540 1878 1717 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03801 1716 1727 1719 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03800 4540 1719 1725 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03799 1725 1727 1723 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03798 1723 1728 1721 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03797 1727 1728 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03796 4540 1726 1728 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03795 1721 1722 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03794 4540 1718 1722 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03793 1878 1716 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03792 4540 1716 1878 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03791 1719 1723 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03790 834 844 836 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03789 4540 877 834 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03788 836 842 835 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03787 4540 835 838 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03786 838 842 837 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03785 837 844 841 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03784 842 844 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03783 4540 839 844 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03782 841 840 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03781 4540 845 840 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03780 877 836 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03779 4540 836 877 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03778 835 837 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03777 214 378 369 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03776 4540 708 214 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03775 369 377 370 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03774 4540 370 217 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03773 217 377 374 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03772 374 378 218 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03771 377 378 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03770 4540 376 378 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03769 218 372 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03768 4540 380 372 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03767 708 369 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03766 4540 369 708 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03765 370 374 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03764 2721 2777 2771 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03763 4540 2802 2721 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03762 2771 2776 2772 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03761 4540 2772 2722 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_03760 2722 2776 2768 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03759 2768 2777 2723 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03758 2776 2777 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03757 4540 2773 2777 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03756 2723 2775 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03755 4540 2774 2775 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03754 2802 2771 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03753 4540 2771 2802 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03752 2772 2768 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_03751 4540 1750 1513 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03750 1513 1894 1600 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03749 1601 2352 1517 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03748 1517 1886 1601 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03747 4540 1600 1517 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03746 1608 1601 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03745 1518 1613 1607 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03744 4540 1886 1518 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03743 1607 1612 1604 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03742 4540 1604 1519 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03741 1519 1612 1606 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03740 1606 1613 1520 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03739 1612 1613 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03738 4540 1609 1613 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03737 1520 1610 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03736 4540 1608 1610 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03735 1886 1607 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03734 4540 1607 1886 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03733 1604 1606 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03732 4540 385 236 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03731 236 537 255 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03730 257 1170 259 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03729 259 1061 257 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03728 4540 255 259 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03727 258 257 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03726 242 250 248 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03725 4540 1061 242 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03724 248 253 247 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03723 4540 247 244 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03722 244 253 245 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03721 245 250 246 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03720 253 250 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03719 4540 249 250 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03718 246 251 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03717 4540 258 251 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03716 1061 248 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03715 4540 248 1061 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03714 247 245 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03713 4540 576 269 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03712 269 855 409 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03711 410 1170 279 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03710 279 1348 410 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03709 4540 409 279 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03708 416 410 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03707 281 422 415 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03706 4540 1348 281 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03705 415 417 412 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03704 4540 412 282 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_03703 282 417 420 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03702 420 422 286 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03701 417 422 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03700 4540 421 422 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03699 286 418 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03698 4540 416 418 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03697 1348 415 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03696 4540 415 1348 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03695 412 420 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_03694 4540 2699 2640 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03693 2640 2655 2641 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03692 2353 2352 2354 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03691 2354 2643 2353 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03690 4540 2641 2354 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03689 2647 2353 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03688 2644 2654 2646 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03687 4540 2643 2644 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03686 2646 2648 2645 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03685 4540 2645 2650 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03684 2650 2648 2651 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03683 2651 2654 2652 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03682 2648 2654 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03681 4540 2653 2654 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03680 2652 2649 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03679 4540 2647 2649 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03678 2643 2646 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03677 4540 2646 2643 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03676 2645 2651 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03675 1733 1894 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03674 1738 1730 1733 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03673 1731 1747 1738 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03672 4540 2315 1731 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03671 1735 1745 1737 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03670 4540 1885 1735 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03669 1737 1743 1736 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03668 4540 1736 1740 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_03667 1740 1743 1741 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03666 1741 1745 1742 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03665 1743 1745 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03664 4540 1744 1745 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03663 1742 1739 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03662 4540 1738 1739 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03661 1885 1737 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03660 4540 1737 1885 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03659 1736 1741 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_03658 538 537 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03657 755 544 538 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03656 540 696 755 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03655 4540 2315 540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03654 525 749 753 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03653 4540 1051 525 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03652 753 748 751 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03651 4540 751 534 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03650 534 748 750 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03649 750 749 532 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03648 748 749 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03647 4540 695 749 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03646 532 758 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03645 4540 755 758 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03644 1051 753 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03643 4540 753 1051 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03642 751 750 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03641 858 855 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03640 867 856 858 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03639 857 859 867 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03638 4540 2315 857 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03637 860 870 861 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03636 4540 1347 860 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03635 861 869 862 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03634 4540 862 863 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03633 863 869 864 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03632 864 870 865 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03631 869 870 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03630 4540 866 870 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03629 865 868 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03628 4540 867 868 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03627 1347 861 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03626 4540 861 1347 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03625 862 864 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03624 2306 2313 2305 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03623 4540 2356 2306 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03622 2305 2309 2303 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03621 4540 2303 2304 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03620 2304 2309 2311 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03619 2311 2313 2310 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03618 2309 2313 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03617 4540 2312 2313 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03616 2310 2308 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03615 4540 2317 2308 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03614 2356 2305 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03613 4540 2305 2356 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03612 2303 2311 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03611 4540 1862 1732 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03610 1732 2002 1863 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03609 1866 2027 1734 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03608 1734 2613 1866 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03607 4540 1863 1734 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03606 1865 1866 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03605 1715 1861 1852 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03604 4540 2027 1715 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03603 1852 1860 1854 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03602 4540 1854 1724 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03601 1724 1860 1857 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03600 1857 1861 1720 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03599 1860 1861 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03598 4540 1859 1861 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03597 1720 1856 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03596 4540 1865 1856 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03595 2027 1852 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03594 4540 1852 2027 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03593 1854 1857 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03592 4540 555 558 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03591 558 765 701 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03590 776 1030 560 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03589 560 2613 776 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03588 4540 701 560 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03587 777 776 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03586 551 767 771 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03585 4540 1030 551 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03584 771 766 769 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03583 4540 769 556 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03582 556 766 768 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03581 768 767 557 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03580 766 767 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03579 4540 700 767 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03578 557 774 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03577 4540 777 774 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03576 1030 771 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03575 4540 771 1030 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03574 769 768 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03573 4540 402 256 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03572 256 853 572 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03571 574 1326 575 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03570 575 2613 574 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03569 4540 572 575 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03568 573 574 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03567 4540 2438 2336 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03566 2336 2497 2333 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03565 2333 2435 2445 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03564 4540 2524 2526 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03563 2441 2450 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03562 2442 2440 2441 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03561 2524 2439 2442 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03560 4540 2438 2344 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03559 2344 2643 2342 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03558 2342 2656 2439 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03557 4540 2438 2340 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03556 2340 2802 2339 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03555 2339 2437 2440 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03554 4540 2198 2073 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03553 2073 2688 2069 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03552 2069 2197 2450 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03551 3111 1355 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03550 1355 1353 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03549 4540 1352 1355 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03548 4540 1368 1264 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03547 1264 1351 1265 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03546 1265 1372 1266 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03545 1266 1350 1353 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03544 4540 1376 1271 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03543 1271 1382 1270 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03542 1270 2696 1368 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03541 4540 1349 1261 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03540 1261 1347 1260 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03539 1260 2357 1351 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03538 4540 1376 1273 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03537 1273 1371 1272 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03536 1272 1911 1372 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03535 4540 1349 1263 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03534 1263 1348 1262 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03533 1262 2656 1350 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03532 4540 1331 1183 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03531 1183 1180 1182 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03530 1182 1214 1181 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03529 1181 1179 1352 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03528 1256 1330 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03527 1254 1441 1331 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03526 1255 1328 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03525 4540 1337 1254 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03524 4540 1326 1253 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03523 1331 2488 1256 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03522 1253 1445 1331 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03521 1331 1329 1255 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03520 1337 1334 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03519 4540 2171 1337 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03518 1445 1442 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03517 4540 2513 1445 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03516 1329 1323 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03515 4540 2325 1329 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03514 1330 1323 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03513 4540 2620 1330 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03512 4540 1152 1143 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03511 1213 1219 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03510 1205 1369 1214 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03509 1210 1206 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03508 4540 1357 1205 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03507 4540 1226 1211 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03506 1214 1232 1213 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03505 1211 1216 1214 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03504 1214 1207 1210 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03503 1369 1376 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03502 4540 2542 1369 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03501 1216 1217 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03500 4540 2220 1216 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03499 1207 1204 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03498 4540 2390 1207 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03497 1219 1217 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03496 4540 2222 1219 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03495 4540 781 1179 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03494 711 709 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03493 712 710 711 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03492 781 713 712 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03491 4540 714 607 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03490 607 723 606 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03489 606 2197 713 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03488 4540 714 588 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03487 588 708 587 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03486 587 1428 710 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03485 4540 714 595 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03484 595 715 596 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03483 596 2447 709 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03482 3377 1060 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03481 1060 1058 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03480 4540 1057 1060 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03479 4540 1070 973 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03478 973 1055 971 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03477 971 1056 972 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03476 972 1066 1058 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03475 4540 1072 983 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03474 983 1091 982 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03473 982 2696 1070 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03472 4540 1166 966 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03471 966 1298 1055 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03470 1166 1164 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03469 4540 2171 1166 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03468 4540 1052 968 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03467 968 1051 967 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03466 967 2357 1056 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03465 4540 930 894 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03464 894 1037 893 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03463 893 898 895 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03462 895 892 1057 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03461 931 929 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03460 925 1377 930 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03459 928 926 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03458 4540 1063 925 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03457 4540 1092 927 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03456 930 1095 931 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03455 927 933 930 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03454 930 1088 928 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03453 1377 1376 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03452 4540 2542 1377 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03451 933 932 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03450 4540 2220 933 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03449 1088 1087 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03448 4540 2390 1088 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03447 929 924 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03446 4540 2222 929 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03445 961 1044 1037 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03444 1037 1032 962 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03443 4540 1030 960 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03442 960 1147 1037 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03441 4540 1033 961 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03440 962 1035 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03439 1147 1145 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03438 4540 2513 1147 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03437 1033 1027 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03436 4540 2325 1033 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03435 1035 1027 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03434 4540 2620 1035 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03433 4540 890 892 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03432 891 888 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03431 889 887 891 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03430 890 1062 889 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03429 3118 2204 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03428 2204 2202 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03427 4540 2203 2204 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03426 2030 2026 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03425 2025 2165 2044 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03424 2029 2027 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03423 4540 2055 2025 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03422 4540 2023 2024 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03421 2044 2168 2030 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03420 2024 2033 2044 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03419 2044 2031 2029 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03418 2165 2166 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03417 4540 2620 2165 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03416 2033 2032 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03415 4540 2171 2033 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03414 4540 2161 2160 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03413 1805 1923 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03412 1800 1920 2042 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03411 1801 2099 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03410 4540 2065 1800 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03409 4540 1915 1802 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03408 2042 1928 1805 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03407 1802 2094 2042 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03406 2042 1914 1801 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03405 4540 2040 2043 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03404 2036 2179 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03403 2039 2035 2036 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03402 2040 2064 2039 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03401 1978 2135 2128 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03400 4540 2516 1978 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03399 2128 2134 2129 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03398 4540 2129 1979 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_03397 1979 2134 2126 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03396 2126 2135 1982 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03395 2134 2135 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03394 4540 2131 2135 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03393 1982 2132 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03392 4540 2130 2132 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03391 2516 2128 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03390 4540 2128 2516 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03389 2129 2126 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_03388 1250 1316 1306 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03387 4540 1328 1250 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03386 1306 1313 1307 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03385 4540 1307 1251 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_03384 1251 1313 1308 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03383 1308 1316 1252 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03382 1313 1316 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03381 4540 1310 1316 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03380 1252 1312 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03379 4540 1311 1312 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03378 1328 1306 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03377 4540 1306 1328 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03376 1307 1308 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_03375 1139 1328 1140 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03374 1140 1585 1139 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03373 4540 1138 1140 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03372 1311 1139 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03371 4540 856 854 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03370 854 853 1138 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03369 202 360 353 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03368 4540 1044 202 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03367 353 362 356 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03366 4540 356 204 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_03365 204 362 358 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03364 358 360 203 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03363 362 360 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03362 4540 359 360 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03361 203 361 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03360 4540 511 361 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03359 1044 353 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03358 4540 353 1044 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03357 356 358 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_03356 4540 513 511 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03355 4540 510 512 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_03354 512 1044 4540 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_03353 513 743 514 4541 tn L=0.32U W=2.45U AS=1.8375P AD=1.8375P PS=6.4U PD=6.4U 
Mtr_03352 514 516 4540 4541 tn L=0.35U W=2.45U AS=1.8865P AD=1.8865P PS=6.45U PD=6.45U 
Mtr_03351 512 745 513 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_03350 1502 1584 1576 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03349 4540 2168 1502 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03348 1576 1583 1575 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03347 4540 1575 1504 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03346 1504 1583 1579 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03345 1579 1584 1505 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03344 1583 1584 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03343 4540 1581 1584 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03342 1505 1577 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03341 4540 1582 1577 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03340 2168 1576 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03339 4540 1576 2168 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03338 1575 1579 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03337 1586 2168 1506 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03336 1506 1585 1586 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03335 4540 1588 1506 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03334 1582 1586 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03333 4540 1730 1508 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03332 1508 2002 1588 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03331 2624 2630 2626 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03330 4540 2636 2624 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03329 2626 2633 2625 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03328 4540 2625 2627 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03327 2627 2633 2628 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03326 2628 2630 2632 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03325 2633 2630 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03324 4540 2629 2630 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03323 2632 2631 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03322 4540 2634 2631 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03321 2636 2626 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03320 4540 2626 2636 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03319 2625 2628 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_03318 2638 2636 2637 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03317 2637 2635 2638 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03316 4540 2639 2637 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03315 2634 2638 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03314 4540 2655 2642 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03313 2642 2841 2639 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03312 1429 1437 1507 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03311 4540 1441 1429 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03310 1507 1436 1509 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03309 4540 1509 1433 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_03308 1433 1436 1510 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03307 1510 1437 1432 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03306 1436 1437 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03305 4540 1434 1437 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03304 1432 1435 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03303 4540 1440 1435 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03302 1441 1507 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03301 4540 1507 1441 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03300 1509 1510 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_03299 4540 1328 1157 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03298 1157 1339 1184 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03297 1184 1156 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03296 1339 1341 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03295 4540 2335 1339 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03294 4540 1154 1156 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03293 1155 2924 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03292 1153 1152 1155 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03291 1154 1159 1153 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03290 4540 1069 981 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03289 981 1067 980 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03288 980 1068 3380 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03287 909 908 912 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03286 4540 907 910 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03285 912 921 911 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03284 910 914 909 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03283 4540 911 1069 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03282 4540 920 906 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03281 906 904 905 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03280 905 1893 907 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03279 4540 920 915 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03278 915 913 916 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03277 916 2934 914 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03276 4540 884 885 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03275 885 1032 886 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03274 886 2812 908 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03273 4540 920 923 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03272 923 926 922 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03271 922 2825 921 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03270 992 1374 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03269 989 1098 1096 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03268 990 1091 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03267 4540 1090 989 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03266 4540 1092 991 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03265 1096 1095 992 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03264 991 1103 1096 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03263 1096 1221 990 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03262 1098 1101 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03261 4540 2229 1098 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03260 1103 1101 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03259 4540 2414 1103 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03258 1221 1222 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03257 4540 1646 1221 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03256 1374 1373 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03255 4540 2410 1374 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03254 4540 707 578 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03253 578 877 577 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03252 577 706 871 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03251 4540 884 876 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03250 876 1030 875 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03249 875 2809 874 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03248 4540 1054 1068 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03247 969 1169 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03246 970 1053 969 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03245 1054 1064 970 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03244 4540 1065 977 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03243 977 1063 976 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03242 976 2814 1064 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03241 964 1051 1053 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03240 1053 1044 965 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03239 4540 1061 963 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03238 963 1338 1053 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03237 4540 1045 964 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03236 965 1049 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03235 1338 1341 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03234 4540 2175 1338 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03233 1045 1042 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03232 4540 1882 1045 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03231 1049 1048 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03230 4540 2335 1049 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03229 4540 1298 1168 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03228 1168 1449 1169 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03227 1169 1167 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03226 1449 1452 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03225 4540 2337 1449 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03224 4540 1163 1167 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03223 1161 2924 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03222 1162 1160 1161 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03221 1163 1159 1162 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03220 4540 2092 2093 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03219 2093 2087 2089 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03218 2089 2088 3221 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03217 4540 2194 2061 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03216 2061 2195 2060 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03215 2060 2827 2196 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03214 4540 2081 2072 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03213 2072 2070 2071 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03212 2071 2934 2076 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03211 4540 2081 2056 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03210 2056 2055 2057 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03209 2057 2812 2075 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03208 4540 2081 2082 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03207 2082 2099 2083 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03206 2083 2825 2084 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03205 1817 1821 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03204 1811 1819 1815 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03203 1814 1812 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03202 4540 1810 1811 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03201 4540 1915 1816 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03200 1815 1928 1817 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03199 1816 1825 1815 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03198 1815 1813 1814 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03197 1819 1824 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03196 4540 2229 1819 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03195 1825 1824 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03194 4540 2414 1825 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03193 1813 1647 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03192 4540 1646 1813 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03191 1821 1824 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03190 4540 2410 1821 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03189 4540 1770 1760 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03188 1760 1878 1759 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03187 1759 2034 1764 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03186 4540 1770 1763 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03185 1763 2027 1761 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03184 1761 2809 1765 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03183 4540 2054 2088 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03182 2051 2170 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03181 2052 2050 2051 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03180 2054 2066 2052 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03179 4540 2081 2067 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03178 2067 2065 2068 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03177 2068 2814 2066 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03176 1767 1886 2050 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03175 2050 2023 1766 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03174 4540 1885 1762 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03173 1762 1884 2050 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03172 4540 1887 1767 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03171 1766 1891 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03170 1884 1881 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03169 4540 1882 1884 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03168 1887 1770 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03167 4540 2175 1887 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03166 1891 1892 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03165 4540 2337 1891 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03164 4540 2168 2028 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03163 2028 2173 2170 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03162 2170 2167 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03161 2173 2172 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03160 4540 2335 2173 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03159 4540 2162 2167 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03158 2018 2924 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03157 2019 2161 2018 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03156 2162 2172 2019 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03155 3289 2669 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03154 2669 2676 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03153 4540 2668 2669 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03152 4540 2671 2673 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03151 2673 2672 2675 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03150 2675 2670 2674 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03149 2674 2680 2676 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03148 4540 2460 2397 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03147 2397 2705 2396 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03146 2396 2696 2671 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03145 4540 2622 2623 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03144 2623 2806 2672 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03143 2622 2621 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03142 4540 2620 2622 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03141 4540 2355 2359 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03140 2359 2356 2358 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03139 2358 2357 2670 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03138 4540 2683 2679 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03137 2679 2677 2678 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03136 2678 2691 2680 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03135 4540 2443 2349 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03134 2349 2444 2351 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03133 2351 2529 2350 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03132 2350 2526 2668 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03131 2389 2388 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03130 2382 2394 2443 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03129 2385 2684 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03128 4540 2664 2382 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03127 4540 2846 2386 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03126 2443 2561 2389 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03125 2386 2384 2443 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03124 2443 2392 2385 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03123 2394 2395 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03122 4540 2542 2394 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03121 2384 2223 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03120 4540 2220 2384 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03119 2392 2391 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03118 4540 2390 2392 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03117 2388 2223 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03116 4540 2222 2388 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03115 2330 2636 2444 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03114 2444 2516 2331 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03113 4540 2801 2326 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03112 2326 2332 2444 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03111 4540 2328 2330 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03110 2331 2327 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03109 2332 2334 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03108 4540 2513 2332 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03107 2328 2166 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03106 4540 2171 2328 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03105 2327 2324 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03104 4540 2325 2327 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03103 4540 2448 2362 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03102 2362 2826 2361 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03101 2361 2447 2449 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03100 4540 1557 1560 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03099 1560 1557 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03098 4540 1559 1557 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03097 1557 3226 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03096 1559 1563 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03095 1558 1563 1557 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03094 1560 1557 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03093 4540 1557 1560 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03092 1563 1561 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03091 4540 1972 1563 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03090 4540 3297 3230 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03089 3230 3297 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03088 4540 3228 3297 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03087 3297 3835 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03086 3228 3232 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03085 3229 3232 3297 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03084 3230 3297 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03083 4540 3297 3230 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03082 3298 3233 3231 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03081 4540 3298 3232 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03080 3231 3299 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03079 4540 2835 2744 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03078 2744 2839 2743 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03077 2743 2834 3560 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03076 2741 2830 2740 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03075 4540 2832 2742 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03074 2740 2831 2833 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03073 2742 2829 2741 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03072 4540 2833 2835 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03071 4540 2828 2739 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03070 2739 2826 2738 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03069 2738 2827 2832 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03068 4540 2687 2690 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03067 2690 2688 2689 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03066 2689 2934 2829 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03065 4540 2807 2735 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03064 2735 2806 2734 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03063 2734 2812 2830 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03062 4540 2687 2686 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03061 2686 2684 2685 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03060 2685 2825 2831 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03059 2838 2837 2745 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03058 4540 2838 2839 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03057 2745 2836 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03056 2408 2411 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03055 2403 2402 2837 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03054 2405 2705 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03053 4540 2677 2403 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03052 4540 2846 2406 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03051 2837 2561 2408 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03050 2406 2416 2837 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03049 2837 2404 2405 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03048 2402 2226 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03047 4540 2229 2402 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03046 2416 2415 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03045 4540 2414 2416 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03044 2404 1647 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03043 4540 1646 2404 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03042 2411 2415 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03041 4540 2410 2411 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03040 2805 2804 2733 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03039 4540 2805 2836 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03038 2733 2803 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03037 4540 2807 2732 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03036 2732 2802 2731 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03035 2731 2811 2804 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03034 4540 2807 2729 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03033 2729 2801 2730 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03032 2730 2809 2803 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03031 4540 2661 2834 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03030 2662 2660 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03029 2663 2659 2662 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03028 2661 2665 2663 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03027 4540 2682 2666 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03026 2666 2664 2667 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03025 2667 2814 2665 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03024 2348 2643 2659 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03023 2659 2636 2347 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03022 4540 2356 2343 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03021 2343 2341 2659 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03020 4540 2345 2348 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03019 2347 2346 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03018 2341 1881 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03017 4540 1882 2341 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03016 2345 2176 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03015 4540 2175 2345 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03014 2346 2338 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03013 4540 2337 2346 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_03012 4540 2516 2329 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03011 2329 2517 2660 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03010 2660 2520 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03009 2517 2338 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03008 4540 2335 2517 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_03007 4540 2519 2520 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03006 2433 2924 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03005 2434 2497 2433 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03004 2519 2436 2434 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_03003 4540 1188 1191 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03002 1191 1193 1190 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03001 1190 1189 3218 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_03000 718 882 717 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02999 4540 716 719 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02998 717 725 782 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02997 719 721 718 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02996 4540 782 1188 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02995 4540 720 610 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02994 610 715 609 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02993 609 1893 716 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02992 4540 720 618 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02991 618 723 619 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02990 619 2934 721 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02989 4540 884 883 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02988 883 2488 881 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02987 881 2812 882 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02986 4540 724 638 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02985 638 1206 639 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02984 639 2825 725 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02983 1234 1396 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02982 1224 1238 1235 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02981 1229 1382 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02980 4540 1371 1224 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02979 4540 1226 1230 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02978 1235 1232 1234 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02977 1230 1231 1235 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02976 1235 1225 1229 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02975 1238 1236 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02974 4540 2229 1238 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02973 1231 1101 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02972 4540 2414 1231 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02971 1225 1222 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02970 4540 1646 1225 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02969 1396 1395 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02968 4540 2410 1396 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02967 4540 707 584 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02966 584 708 585 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02965 585 706 1175 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02964 4540 1172 1174 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02963 1174 1326 1173 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02962 1173 2809 1176 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02961 4540 1187 1189 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02960 1185 1184 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02959 1186 1345 1185 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02958 1187 1196 1186 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02957 4540 1198 1199 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02956 1199 1357 1195 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02955 1195 2814 1196 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02954 1257 1348 1345 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02953 1345 1441 1259 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02952 4540 1347 1258 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02951 1258 1451 1345 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02950 4540 1343 1257 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02949 1259 1454 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02948 1451 1452 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02947 4540 1882 1451 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02946 1343 1341 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02945 4540 2175 1343 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02944 1454 1452 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02943 4540 2337 1454 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02942 3800 3798 3801 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02941 4540 3800 3797 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02940 3801 3808 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02939 4540 4041 4043 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02938 4043 4329 4044 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02937 4540 4122 4074 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02936 4074 4123 4073 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02935 4073 4343 4221 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02934 4540 4119 4120 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02933 4120 4214 4123 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02932 4344 4345 4346 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02931 4346 4342 4344 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02930 4344 4341 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02929 4333 4331 4330 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02928 4540 4333 4338 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02927 4330 4347 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02926 4058 3912 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02925 3912 3915 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02924 4540 3914 3912 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02923 4540 4070 4066 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02922 4067 4066 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02921 4540 4214 4067 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02920 4337 3803 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02919 3803 3802 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02918 4540 3916 3803 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02917 4540 3915 3916 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02916 4540 4117 4345 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02915 4540 4337 4341 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02914 4540 4058 3917 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02913 3804 3808 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02912 4540 3916 3804 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02911 4065 4064 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02910 4064 4337 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02909 4540 4067 4064 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02908 4061 4059 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02907 4061 4058 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02906 4540 4067 4061 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02905 4540 4061 4122 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02904 4059 3226 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02903 4540 3299 4059 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02902 4053 3905 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02901 4540 3908 4053 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02900 4055 4053 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02899 4055 4058 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02898 4540 4338 4055 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02897 4540 4055 4054 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02896 4540 4054 4046 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02895 4046 4044 4047 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02894 4047 4051 4210 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02893 4339 4340 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02892 4340 4337 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02891 4540 4338 4340 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02890 4056 3908 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02889 4540 3911 4056 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02888 4540 4324 4328 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02887 4328 4325 4326 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02886 4326 4332 4327 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02885 3805 3808 3806 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02884 3806 3835 3805 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02883 3805 3917 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02882 4072 4071 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02881 4540 4070 4072 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02880 4540 4068 3815 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02879 3815 3813 3816 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02878 3816 3814 3921 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02877 4051 4049 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02876 4540 4065 4049 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02875 4052 4320 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02874 4049 4345 4052 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02873 4343 4349 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02872 4540 4346 4349 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02871 4348 4347 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02870 4349 4345 4348 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02869 4332 4336 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02868 4540 4339 4336 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02867 4335 4334 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02866 4336 4345 4335 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02865 4540 4321 4323 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02864 4323 4322 4325 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02863 4057 4056 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02862 4057 4058 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02861 4540 4213 4057 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02860 4540 4057 4324 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02859 4540 3659 3571 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02858 3571 3918 3813 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02857 4069 4072 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02856 4069 4337 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02855 4540 4213 4069 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02854 4540 4069 4068 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02853 3814 3809 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02852 4540 3806 3809 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02851 3812 4334 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02850 3809 3808 3812 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02849 4212 4117 4116 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02848 4540 4212 4213 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02847 4116 4320 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02846 4540 3918 4334 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02845 4540 4322 4320 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02844 4540 4329 4347 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02843 4540 3652 3931 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02842 3931 3652 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02841 4540 3653 3652 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02840 3652 4214 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02839 3653 3804 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02838 3654 3804 3652 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02837 3931 3652 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02836 4540 3652 3931 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02835 4540 3796 4084 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02834 4084 3796 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02833 4540 3794 3796 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02832 3796 3918 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02831 3794 3797 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02830 3795 3797 3796 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02829 4084 3796 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02828 4540 3796 4084 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02827 4540 3790 3792 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02826 3790 3918 4540 4541 tn L=0.35U W=0.75U AS=0.5775P AD=0.5775P PS=3.05U PD=3.05U 
Mtr_02825 4540 3903 3904 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02824 3903 4322 4540 4541 tn L=0.32U W=0.75U AS=0.5625P AD=0.5625P PS=3U PD=3U 
Mtr_02823 4540 3910 3907 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02822 3910 4329 4540 4541 tn L=0.32U W=0.75U AS=0.5625P AD=0.5625P PS=3U PD=3U 
Mtr_02821 4060 4216 4220 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02820 4540 4214 4060 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02819 4220 4215 4219 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02818 4540 4219 4062 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_02817 4062 4215 4217 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02816 4217 4216 4063 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02815 4215 4216 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02814 4540 4118 4216 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02813 4063 4224 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02812 4540 4221 4224 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02811 4214 4220 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02810 4540 4220 4214 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02809 4219 4217 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_02808 4045 4203 4205 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02807 4540 4329 4045 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02806 4205 4202 4208 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02805 4540 4208 4050 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_02804 4050 4202 4206 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02803 4206 4203 4048 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02802 4202 4203 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02801 4540 4115 4203 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02800 4048 4211 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02799 4540 4210 4211 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02798 4329 4205 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02797 4540 4205 4329 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02796 4208 4206 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_02795 4310 4317 4311 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02794 4540 4322 4310 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02793 4311 4319 4312 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02792 4540 4312 4314 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_02791 4314 4319 4313 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02790 4313 4317 4315 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02789 4319 4317 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02788 4540 4316 4317 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02787 4315 4318 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02786 4540 4327 4318 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02785 4322 4311 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02784 4540 4311 4322 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02783 4312 4313 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_02782 3807 3928 3920 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02781 4540 3918 3807 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02780 3920 3929 3922 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02779 4540 3922 3810 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_02778 3810 3929 3925 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02777 3925 3928 3811 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02776 3929 3928 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02775 4540 3926 3928 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02774 3811 3927 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02773 4540 3921 3927 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02772 3918 3920 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02771 4540 3920 3918 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02770 3922 3925 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_02769 4540 3656 3655 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02768 3656 4214 4540 4541 tn L=0.32U W=0.75U AS=0.5625P AD=0.5625P PS=3U PD=3U 
Mtr_02767 4540 3045 3044 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02766 4540 3902 3880 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02765 4540 3209 3269 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02764 4540 3521 3246 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02763 3246 4107 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02762 3319 3479 3246 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02761 3246 4232 3319 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02760 4540 3521 3248 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02759 3248 4232 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02758 3322 3599 3248 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02757 3248 4107 3322 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02756 4540 3073 3254 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02755 4540 3367 3103 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02754 4540 4292 4293 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02753 4540 2786 4269 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02752 3734 3852 3732 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02751 3732 3729 3734 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02750 3734 3983 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02749 4540 3726 3725 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02748 3725 3844 3722 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02747 3722 3732 3723 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02746 3723 3733 3724 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02745 4540 4259 4260 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02744 4540 4161 4009 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02743 4009 4279 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02742 4164 4163 4009 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02741 4009 4269 4164 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02740 4540 3694 3587 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02739 3871 3869 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02738 3869 4167 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02737 4540 4016 3869 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02736 4540 3760 3522 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02735 3522 3520 3521 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02734 3521 3515 3519 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02733 3519 3516 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02732 4540 3516 3520 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02731 3515 3760 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02730 3762 4283 3761 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02729 4540 3766 3763 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02728 3761 3771 3764 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02727 3763 3772 3762 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02726 4540 3764 3760 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02725 4540 4196 3767 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02724 3767 4163 3765 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02723 3765 4187 3766 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02722 4540 3886 3773 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02721 3773 4287 3772 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02720 4540 3774 3770 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02719 3770 4105 3771 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02718 2898 2897 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02717 2897 2916 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02716 4540 3431 2897 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02715 3045 3032 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02714 3032 3031 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02713 4540 4233 3032 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02712 2876 2875 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02711 2875 2873 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02710 4540 4137 2875 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02709 4008 4007 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02708 4007 4186 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02707 4540 4010 4007 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02706 4540 4261 4087 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02705 4087 4269 4090 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02704 4540 4261 4004 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02703 4004 4104 4005 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02702 4540 4241 4240 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02701 4540 4096 4261 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02700 3580 3584 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02699 4540 4232 3579 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02698 3462 3579 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02697 3578 3580 3462 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02696 3465 4232 3578 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02695 4540 3584 3465 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02694 4195 4198 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02693 4540 4196 4194 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02692 4040 4194 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02691 4308 4195 4040 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02690 4042 4196 4308 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02689 4540 4198 4042 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02688 4309 4308 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02687 4540 4303 4307 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02686 4304 4307 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02685 4305 4309 4304 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02684 4306 4303 4305 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02683 4540 4308 4306 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02682 4189 4198 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02681 4540 4196 4190 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02680 4031 4190 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02679 4191 4189 4031 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02678 4036 4196 4191 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02677 4540 4198 4036 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02676 4037 4032 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02675 4540 4191 4030 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02674 4033 4030 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02673 4034 4037 4033 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02672 4035 4191 4034 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02671 4540 4032 4035 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02670 3283 3635 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02669 4540 3638 3282 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02668 3213 3282 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02667 3277 3283 3213 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02666 3212 3638 3277 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02665 4540 3635 3212 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02664 3275 3277 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02663 4540 3276 3278 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02662 3208 3278 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02661 3209 3275 3208 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02660 3210 3276 3209 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02659 4540 3277 3210 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02658 4540 3532 3075 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02657 3078 3075 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02656 4540 3431 3078 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02655 3778 3886 3779 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02654 4540 3778 3774 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02653 3779 4298 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02652 4540 4016 3886 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02651 3839 2883 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02650 2883 2881 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02649 4540 3503 2883 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02648 3698 4137 3699 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02647 4540 3698 3840 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02646 3699 4107 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02645 4137 3071 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02644 3071 3070 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02643 4540 3781 3071 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02642 3787 3786 3788 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02641 4540 3787 3785 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02640 3788 4187 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02639 3783 3786 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02638 4540 4187 3783 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02637 3783 4039 3782 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02636 3782 3785 3783 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02635 4540 3782 3781 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02634 4540 4144 3994 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02633 4233 3998 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02632 3998 4010 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02631 4540 4024 3998 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02630 4029 4198 4027 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02629 4540 4029 4028 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02628 4027 4303 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02627 4026 4303 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02626 4540 4198 4026 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02625 4026 4039 4025 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02624 4025 4028 4026 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02623 4540 4025 4024 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02622 3348 3619 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02621 4540 3367 3348 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02620 4540 3345 3348 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02619 3348 3344 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02618 3506 3348 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02617 3434 3623 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02616 4540 4269 3434 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02615 3434 3514 3505 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02614 3505 3506 3434 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02613 4540 3505 3614 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02612 3343 3342 3256 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02611 4540 3343 3345 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02610 3256 3353 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02609 3623 3356 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02608 3356 3537 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02607 4540 3355 3356 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02606 4540 4258 4262 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02605 3499 2895 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02604 2895 2916 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02603 4540 3070 2895 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02602 2915 3786 2914 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02601 4540 2915 2916 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02600 2914 3103 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02599 4540 3509 3882 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02598 4540 3110 3537 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02597 3510 3537 3513 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02596 4540 3510 3514 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02595 3513 3882 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02594 4540 3710 3500 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02593 3500 3712 3619 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02592 4540 3532 3786 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02591 3353 3786 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02590 4540 3509 3353 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02589 4540 3492 3592 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02588 3255 3181 3176 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02587 4540 3255 3583 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02586 3176 3492 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02585 3181 4269 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02584 4540 4232 3181 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02583 4540 3514 3181 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02582 3181 3355 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02581 4540 3829 3503 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02580 4540 3714 4163 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02579 4540 4301 4302 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02578 4540 4298 4303 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02577 4300 4302 4299 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02576 4540 4300 4297 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02575 4299 4298 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02574 4172 4297 4106 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02573 4540 4172 4272 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02572 4106 4105 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02571 4540 4032 4287 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02570 4540 4289 4285 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02569 4540 4284 4273 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02568 4540 3727 4283 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02567 4540 4283 4110 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02566 4110 4273 4177 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02565 4286 4284 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02564 4286 4285 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02563 4540 4283 4286 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02562 4540 4286 4295 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02561 4015 4273 4014 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02560 4540 4015 4280 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02559 4014 4032 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02558 4281 4290 4282 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02557 4540 4281 4279 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02556 4282 4280 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02555 4185 4303 4114 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02554 4540 4185 4186 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02553 4114 4273 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02552 4540 4104 4167 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02551 4011 4163 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02550 4540 4301 4011 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02549 4540 4186 4011 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02548 4011 4167 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02547 4161 4011 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02546 4019 4287 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02545 4540 4187 4019 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02544 4019 4196 4018 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02543 4018 4020 4019 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02542 4540 4018 4146 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02541 4022 4287 4021 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02540 4540 4022 4020 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02539 4021 4187 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02538 4148 4272 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02537 4540 4146 4148 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02536 3694 3696 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02535 3696 3690 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02534 4540 3983 3696 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02533 3440 3537 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02532 4540 4198 3440 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02531 3440 4196 3525 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02530 3525 3531 3440 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02529 4540 3525 3526 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02528 3529 4198 3530 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02527 4540 3529 3531 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02526 3530 3537 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02525 4540 3331 3325 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02524 3597 3727 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02523 4540 3594 3596 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02522 3485 3596 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02521 3599 3597 3485 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02520 3484 3594 3599 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02519 4540 3727 3484 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02518 4540 4179 4023 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02517 4023 4180 4182 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02516 4182 4296 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02515 4540 4293 4296 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02514 4296 4294 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02513 4296 4295 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02512 4013 4280 4012 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02511 4540 4013 4010 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02510 4012 4105 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02509 2918 3103 2917 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02508 4540 2918 2919 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02507 2917 3110 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02506 4540 2800 3070 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02505 4540 4038 4105 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02504 4540 3502 3846 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02503 4540 2886 4243 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02502 4540 4232 4107 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02501 4540 4198 4187 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02500 4540 3638 3636 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02499 4540 3991 3983 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02498 4540 4196 4039 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02497 4540 3635 3637 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02496 4259 4285 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02495 4540 4272 4259 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02494 4278 4262 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02493 4540 4261 4278 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02492 4540 3171 3160 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02491 3160 4107 3310 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02490 4258 4253 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02489 4540 4252 4258 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02488 4104 4102 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02487 4540 3999 4104 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02486 4241 4253 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02485 4540 4261 4241 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02484 4540 3710 3706 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02483 3706 3705 4096 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02482 4096 3709 3704 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02481 3704 3712 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02480 4540 3712 3705 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02479 3709 3710 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02478 4540 4233 3141 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02477 3141 4269 3239 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02476 2867 4137 2866 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02475 4540 2867 2868 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02474 2866 4269 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02473 4540 4198 3791 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02472 3791 3899 3902 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02471 3902 3900 3789 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02470 3789 4196 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02469 4540 4196 3899 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02468 3900 4198 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02467 4540 4105 2999 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02466 2999 3078 3073 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02465 3073 3077 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02464 4540 4163 4017 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02463 4017 4302 4016 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02462 4540 3882 3430 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02461 3430 3503 3431 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02460 3584 3594 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02459 4540 4148 3584 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02458 4540 3353 3182 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02457 3182 4105 3492 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02456 3331 3619 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02455 4540 4269 3331 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02454 3747 3745 3746 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02453 4540 3747 3744 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02452 3746 4283 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02451 3864 3862 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02450 3862 3871 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02449 4540 4280 3862 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02448 3742 3741 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02447 3741 4280 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02446 4540 4269 3741 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02445 3192 3189 3262 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02444 4540 3846 3192 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02443 3191 3190 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02442 3262 3625 3191 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02441 4540 3262 3188 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02440 4540 3083 3001 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02439 3001 3082 3000 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02438 3000 3098 3189 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02437 3081 3078 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02436 3081 3077 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02435 4540 3091 3081 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02434 4540 3081 3083 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02433 4540 3983 2892 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02432 2892 4269 2891 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02431 2891 2890 3082 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02430 4540 4232 2889 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02429 2889 2885 2890 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02428 2890 2888 2884 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02427 2884 2886 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02426 4540 2886 2885 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02425 2888 4232 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02424 3102 4243 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02423 3102 3096 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02422 4540 3774 3102 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02421 4540 3102 3098 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02420 4540 3624 3523 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02419 3523 4111 3524 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02418 3524 3630 3625 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02417 4540 3626 3517 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02416 3517 3633 3518 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02415 3518 3623 3624 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02414 4113 4179 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_02413 4112 4243 4111 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02412 4540 4113 4112 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02411 3533 3634 3630 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02410 3630 3629 3533 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02409 3533 3991 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02408 3634 4102 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02407 4540 3633 3634 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02406 4540 3628 3629 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02405 3528 3633 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02404 3527 4102 3528 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02403 3628 3627 3527 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02402 4540 4232 4095 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02401 4095 4233 4098 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02400 4144 4143 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02399 4540 4163 4144 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02398 4540 3710 3711 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02397 3714 3711 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02396 4540 3712 3714 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02395 4540 2919 2728 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02394 2728 4105 2800 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02393 3829 3710 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02392 4540 3712 3829 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02391 4179 4177 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02390 4540 4287 4179 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02389 4540 4290 4291 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02388 4291 4297 4292 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02387 4540 3638 3541 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02386 3541 3637 4298 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02385 4540 4287 4288 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02384 4288 4302 4289 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02383 4301 4196 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02382 4540 4187 4301 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02381 4540 3635 3540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02380 3540 3636 4032 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02379 4284 4198 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02378 4540 4039 4284 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02377 4540 3712 3601 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02376 3727 3601 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02375 4540 3710 3727 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02374 4540 3619 3002 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02373 3002 3103 3355 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02372 4540 3636 3442 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02371 3442 3637 3532 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02370 3509 4198 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02369 4540 4196 3509 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02368 4540 3638 2935 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02367 2935 3635 3110 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02366 3366 4198 3267 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02365 4540 3366 3367 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02364 3267 4196 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02363 2790 3835 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02362 4540 3226 2790 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02361 4540 3905 2790 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02360 2790 3911 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02359 4540 3657 3658 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02358 3657 3835 4540 4541 tn L=0.35U W=0.75U AS=0.5775P AD=0.5775P PS=3.05U PD=3.05U 
Mtr_02357 3743 4182 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02356 4540 4107 3743 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02355 3743 4010 3868 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02354 3868 4161 3743 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02353 4540 3868 3865 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02352 3737 4269 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02351 4540 3735 3737 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02350 3737 4243 3736 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02349 3736 3865 3737 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02348 4540 3736 3733 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02347 3621 4167 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02346 4540 3619 3621 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02345 3616 3614 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02344 4540 4107 3616 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02343 3617 3616 3508 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02342 3508 3621 3617 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02341 4540 4243 3508 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02340 3729 3617 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02339 4001 4102 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02338 4540 4182 4001 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02337 4263 4262 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02336 4540 4283 4263 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02335 3854 4263 3728 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02334 3728 4001 3854 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02333 4540 3850 3728 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02332 3852 3854 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02331 4540 4141 4142 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02330 4099 4144 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02329 4100 4098 4099 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02328 4141 4101 4100 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02327 4540 3840 3843 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02326 3843 3850 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02325 3843 3839 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02324 3713 3843 3844 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02323 3844 4142 3713 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02322 3713 3991 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02321 3606 4262 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02320 4540 3509 3606 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02319 4540 3503 3606 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02318 3606 3499 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02317 3608 4102 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02316 4540 3614 3608 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02315 3497 3608 3726 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02314 3726 3606 3497 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02313 3497 4243 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02312 4540 4272 4264 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02311 4264 4294 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02310 4264 4295 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02309 4540 4260 4157 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02308 4157 4269 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02307 4157 4177 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02306 4154 4157 4002 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02305 4002 4264 4154 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02304 4540 4102 4002 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02303 4152 4154 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02302 4000 4164 4150 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02301 4150 4152 4000 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02300 4000 4243 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02299 3326 3327 3250 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02298 4540 3326 3486 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02297 3250 3325 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02296 4540 4269 3489 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02295 3489 3526 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02294 3489 3592 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02293 3487 3489 3419 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02292 3419 4107 3487 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02291 4540 3486 3419 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02290 3488 3487 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02289 3468 3466 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02288 3466 4232 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02287 4540 4148 3466 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02286 4540 3467 3470 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02285 3411 3468 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02284 3412 3599 3411 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02283 3467 4243 3412 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02282 3474 3470 3701 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02281 3701 3488 3474 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02280 3474 3983 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02279 3595 3594 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02278 4540 3592 3595 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02277 3585 3584 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_02276 3469 4232 3591 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02275 4540 3585 3469 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02274 4540 3583 3473 4541 tn L=0.35U W=2.45U AS=1.8865P AD=1.8865P PS=6.45U PD=6.45U 
Mtr_02273 3473 3829 4540 4541 tn L=0.35U W=2.45U AS=1.8865P AD=1.8865P PS=6.45U PD=6.45U 
Mtr_02272 4540 3595 3473 4541 tn L=0.32U W=2.45U AS=1.8375P AD=1.8375P PS=6.4U PD=6.4U 
Mtr_02271 3473 3586 3700 4541 tn L=0.32U W=2.45U AS=1.8375P AD=1.8375P PS=6.4U PD=6.4U 
Mtr_02270 3700 3714 3471 4541 tn L=0.32U W=3.32U AS=2.49P AD=2.49P PS=8.15U PD=8.15U 
Mtr_02269 3471 3587 3472 4541 tn L=0.35U W=3.32U AS=2.5564P AD=2.5564P PS=8.2U PD=8.2U 
Mtr_02268 3472 3591 4540 4541 tn L=0.32U W=3.32U AS=2.49P AD=2.49P PS=8.15U PD=8.15U 
Mtr_02267 4540 3700 3703 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02266 3703 3701 3702 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02265 3702 4150 3716 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02264 3721 3716 3720 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02263 4540 3717 3721 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02262 3719 3846 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02261 3720 3724 3719 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02260 4540 3720 3715 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02259 4540 2868 2869 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02258 4540 3239 3038 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02257 4540 4243 3754 4541 tn L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mtr_02256 3749 3846 4540 4541 tn L=0.32U W=0.72U AS=0.54P AD=0.54P PS=2.95U PD=2.95U 
Mtr_02255 3759 3748 3753 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02254 3753 4243 3752 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02253 3752 3754 3758 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02252 3758 3887 3759 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02251 4540 3846 3759 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02250 3751 3749 4540 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02249 3752 3872 3751 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02248 4540 3752 3905 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02247 4540 4269 3875 4541 tn L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mtr_02246 3874 4243 4540 4541 tn L=0.32U W=0.72U AS=0.54P AD=0.54P PS=2.95U PD=2.95U 
Mtr_02245 3757 3896 3755 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02244 3755 4269 3877 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02243 3877 3875 3756 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02242 3756 3880 3757 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02241 4540 4243 3757 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02240 3750 3874 4540 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02239 3877 3881 3750 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02238 4540 3877 3872 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02237 3769 3902 3883 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02236 4540 3884 3769 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02235 3768 4269 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02234 3883 3882 3768 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02233 4540 3883 3881 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02232 4540 4305 3784 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02231 3784 3895 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02230 3896 4034 3784 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02229 3784 4105 3896 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02228 4540 3362 3363 4541 tn L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mtr_02227 3358 4269 4540 4541 tn L=0.32U W=0.72U AS=0.54P AD=0.54P PS=2.95U PD=2.95U 
Mtr_02226 3266 3370 3264 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02225 3264 3362 3360 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02224 3360 3363 3265 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02223 3265 3538 3266 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02222 4540 4269 3266 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02221 3263 3358 4540 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02220 3360 3367 3263 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02219 4540 3360 3748 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02218 3369 3532 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02217 4540 3372 3368 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02216 3271 3368 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02215 3370 3369 3271 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02214 3273 3372 3370 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02213 4540 3532 3273 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02212 3375 4198 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02211 4540 4196 3373 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02210 3274 3373 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02209 3372 3375 3274 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02208 3279 4196 3372 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02207 4540 4198 3279 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02206 3535 3548 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02205 4540 3537 3534 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02204 3536 3534 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02203 3538 3535 3536 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02202 3539 3537 3538 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02201 4540 3548 3539 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02200 3543 4198 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02199 4540 4196 3542 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02198 3546 3542 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02197 3548 3543 3546 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02196 3549 4196 3548 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02195 4540 4198 3549 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02194 4540 4105 3893 4541 tn L=0.35U W=1.02U AS=0.7854P AD=0.7854P PS=3.6U PD=3.6U 
Mtr_02193 3888 4269 4540 4541 tn L=0.35U W=0.72U AS=0.5544P AD=0.5544P PS=3U PD=3U 
Mtr_02192 3780 4034 3776 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_02191 3776 4105 3891 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_02190 3891 3893 3777 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_02189 3777 4305 3780 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_02188 4540 4269 3780 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_02187 3775 3888 4540 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_02186 3891 4284 3775 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_02185 4540 3891 3887 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02184 4540 3091 3087 4541 tn L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mtr_02183 3086 3084 4540 4541 tn L=0.32U W=0.72U AS=0.54P AD=0.54P PS=2.95U PD=2.95U 
Mtr_02182 3006 3085 3004 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02181 3004 3091 3089 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02180 3089 3087 3005 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02179 3005 3109 3006 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02178 4540 3084 3006 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02177 3003 3086 4540 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02176 3089 3194 3003 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02175 4540 3089 3226 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02174 4540 4269 3201 4541 tn L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mtr_02173 3195 4243 4540 4541 tn L=0.32U W=0.72U AS=0.54P AD=0.54P PS=2.95U PD=2.95U 
Mtr_02172 3202 3209 3198 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02171 3198 4269 3197 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02170 3197 3201 3199 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02169 3199 3537 3202 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02168 4540 4243 3202 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02167 3196 3195 4540 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02166 3197 3200 3196 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02165 4540 3197 3194 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02164 4540 4287 3205 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_02163 3205 3272 3270 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_02162 4540 3272 3268 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_02161 3270 3268 3206 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_02160 3206 3269 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_02159 3200 3270 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02158 4540 3786 2923 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02157 2923 2926 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02156 3085 2944 2923 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02155 2923 4269 3085 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02154 2946 3638 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02153 4540 3635 2943 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02152 2942 2943 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02151 2944 2946 2942 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02150 2947 3635 2944 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02149 4540 3638 2947 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02148 4540 3106 3008 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02147 3008 3104 3109 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02146 3109 3107 3007 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02145 3007 3105 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02144 4540 3105 3104 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02143 3107 3106 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02142 2941 3635 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02141 4540 3638 2938 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02140 2936 2938 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02139 3106 2941 2936 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02138 2940 3638 3106 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02137 4540 3635 2940 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02136 3105 2928 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02135 2928 2925 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02134 4540 2926 2928 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02133 4540 3991 3057 4541 tn L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mtr_02132 3056 3055 4540 4541 tn L=0.32U W=0.72U AS=0.54P AD=0.54P PS=2.95U PD=2.95U 
Mtr_02131 2993 3158 2994 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02130 2994 3991 3059 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02129 3059 3057 2992 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02128 2992 3165 2993 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02127 4540 3055 2993 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02126 2991 3056 4540 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02125 3059 3065 2991 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02124 4540 3059 4397 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02123 3065 3069 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02122 4540 3064 2996 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02121 2996 3991 3069 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02120 2997 4243 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02119 4540 3091 2998 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02118 3069 3066 2997 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02117 2998 3855 3069 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02116 4540 3052 2990 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02115 2990 3053 3064 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02114 4540 3049 2989 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02113 2989 3994 2988 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02112 2988 3048 3052 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02111 4540 4232 2987 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02110 2987 3045 3048 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02109 4540 4243 2880 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02108 2880 3839 2879 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02107 2879 2878 3053 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02106 4540 2876 2877 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02105 2877 4107 2878 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02104 4540 4283 3730 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02103 3730 3861 3731 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02102 3731 3858 3855 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02101 3861 3859 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02100 3859 4008 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02099 4540 3871 3859 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02098 3858 3856 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02097 3856 4010 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02096 4540 4269 3856 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02095 4540 3619 2726 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02094 2726 2792 2725 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02093 2725 2798 3066 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02092 2794 2898 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02091 2794 3253 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02090 4540 3070 2794 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02089 4540 2794 2792 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02088 4540 2799 2727 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02087 2727 2800 2798 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02086 3158 3247 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02085 4540 3164 3247 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02084 3159 3319 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02083 3247 4243 3159 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02082 4540 3714 3480 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02081 3480 3475 3479 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02080 3479 3476 3478 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02079 3478 3477 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02078 4540 3477 3475 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02077 3476 3714 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02076 4540 4243 3164 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02075 3164 3583 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02074 3164 3161 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02073 4540 3503 2995 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02072 2995 3062 3161 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02071 3161 3073 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02070 4540 3169 3165 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02069 4540 3174 3170 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_02068 3170 3177 4540 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_02067 3169 4243 3168 4541 tn L=0.35U W=2.45U AS=1.8865P AD=1.8865P PS=6.45U PD=6.45U 
Mtr_02066 3168 3322 4540 4541 tn L=0.32U W=2.45U AS=1.8375P AD=1.8375P PS=6.4U PD=6.4U 
Mtr_02065 3170 3172 3169 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_02064 4540 4167 3175 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02063 3175 3325 3173 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02062 3173 3254 3174 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02061 3177 4269 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02060 4540 4107 3177 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02059 4540 2898 3177 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02058 3177 2900 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02057 2901 2925 2899 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02056 4540 2901 2900 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02055 2899 2919 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02054 3493 3498 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02053 3426 3613 3498 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_02052 4540 3495 3426 4541 tn L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mtr_02051 3426 3847 4540 4541 tn L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mtr_02050 4540 3983 3426 4541 tn L=0.32U W=1.02U AS=0.765P AD=0.765P PS=3.55U PD=3.55U 
Mtr_02049 3498 3603 3424 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mtr_02048 3424 3502 3425 4541 tn L=0.35U W=2.17U AS=1.6709P AD=1.6709P PS=5.9U PD=5.9U 
Mtr_02047 3425 3496 4540 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mtr_02046 4540 3622 3435 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02045 3435 3507 3496 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02044 4540 4243 3511 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02043 3511 4163 3512 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02042 3512 4174 3622 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02041 4173 4107 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02040 4173 4177 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02039 4540 4297 4173 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02038 4540 4173 4174 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02037 4540 3260 3186 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02036 3186 3352 3185 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02035 3185 3258 3507 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02034 3260 3261 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02033 3261 3272 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02032 4540 3353 3261 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02031 3351 3350 3259 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02030 4540 3351 3352 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02029 3259 3503 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02028 3257 3355 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02027 3257 3310 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02026 4540 3353 3257 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_02025 4540 3257 3258 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02024 4540 3983 3490 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02023 3490 3602 3491 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02022 3491 3604 3603 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02021 3251 3329 3602 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02020 3602 3331 3251 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02019 3251 3327 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02018 4540 3781 3252 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02017 3252 3344 3329 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02016 3329 4107 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02015 3494 3851 3604 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02014 3604 3727 3494 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02013 3494 4243 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02012 3851 4102 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02011 4540 4024 3851 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02010 4540 3481 3483 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02009 3483 3839 3495 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02008 3495 3482 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02007 3481 3323 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_02006 4540 4232 3323 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02005 3249 4269 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02004 3323 3526 3249 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_02003 4540 3996 3718 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02002 3718 3994 3847 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02001 3847 4243 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_02000 3996 3997 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01999 4540 4252 3997 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01998 3995 4269 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01997 3997 4146 3995 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01996 4540 3611 3504 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01995 3504 3740 3613 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01994 3613 3610 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01993 4540 2913 2908 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01992 2908 2907 2906 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01991 2906 2905 3611 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01990 2912 3619 2911 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01989 4540 2912 2913 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01988 2911 4243 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01987 2907 2910 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01986 2910 2919 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01985 4540 4269 2910 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01984 2904 3431 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01983 2904 3253 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01982 4540 2919 2904 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01981 4540 2904 2905 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01980 4540 3744 3738 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01979 3738 3864 3739 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01978 3739 3742 3740 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01977 4540 3837 3835 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01976 4540 4246 3708 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_01975 3708 3833 4540 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_01974 3837 3846 3707 4541 tn L=0.32U W=2.45U AS=1.8375P AD=1.8375P PS=6.4U PD=6.4U 
Mtr_01973 3707 3981 4540 4541 tn L=0.35U W=2.45U AS=1.8865P AD=1.8865P PS=6.45U PD=6.45U 
Mtr_01972 3708 3836 3837 4541 tn L=0.32U W=1.6U AS=1.2P AD=1.2P PS=4.7U PD=4.7U 
Mtr_01971 3987 3986 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01970 4540 3982 3984 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01969 3985 4092 3988 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01968 4540 3983 3985 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01967 3981 3988 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01966 3988 4243 3987 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01965 3984 3991 3988 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01964 3988 4265 3989 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01963 3989 3990 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01962 4540 4238 4093 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01961 4093 4135 4092 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01960 4540 4235 4239 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01959 4239 4241 4237 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01958 4237 4236 4238 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01957 4236 4234 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01956 4234 4232 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01955 4540 4233 4234 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01954 4134 4139 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01953 4134 4088 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01952 4540 4090 4134 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01951 4540 4134 4135 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01950 4139 4137 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01949 4540 4252 4139 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01948 4540 3973 3975 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01947 3975 4132 3982 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01946 3820 4240 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01945 3820 3840 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01944 4540 3819 3820 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01943 4540 3820 3973 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01942 4131 4094 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01941 4131 4243 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01940 4540 4090 4131 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01939 4540 4131 4132 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01938 4540 4098 4094 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01937 3334 3336 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01936 3334 3331 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01935 4540 3341 3334 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01934 4540 3334 3986 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01933 3341 3345 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01932 4540 3367 3341 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01931 4540 4005 3341 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01930 3341 3514 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01929 4540 3509 3336 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01928 3336 3499 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01927 3336 4003 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01926 4540 4278 4003 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01925 4540 4270 4267 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01924 4267 4275 4268 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01923 4268 4266 4265 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01922 4270 4271 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01921 4271 4283 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01920 4540 4269 4271 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01919 4540 4278 4277 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01918 4277 4292 4276 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01917 4276 4273 4274 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01916 4274 4289 4275 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01915 4006 4301 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01914 4006 4008 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01913 4540 4005 4006 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01912 4540 4006 4266 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01911 4245 4250 4244 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01910 4540 4245 4246 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01909 4244 4243 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01908 4540 4247 4251 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01907 4251 4256 4249 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01906 4249 4248 4250 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01905 4540 4253 4242 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01904 4242 4261 4247 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01903 4540 4273 4257 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01902 4257 4259 4254 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01901 4254 4261 4255 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01900 4255 4258 4256 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01899 4540 4096 4097 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01898 4097 4169 4248 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01897 4169 4186 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01896 4540 4279 4169 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01895 4540 4301 4169 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01894 4169 4167 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01893 4540 3823 3695 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01892 3695 3972 3693 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01891 3693 3824 3833 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01890 3692 3691 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01889 3692 3694 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01888 4540 4240 3692 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01887 4540 3692 3823 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01886 3689 4232 3688 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01885 4540 3689 3691 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01884 3688 4148 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01883 3974 4232 3972 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01882 3972 3977 3974 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01881 3974 3980 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01880 3979 4148 3976 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01879 4540 3979 3977 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01878 3976 4269 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01877 4540 4261 3978 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01876 3980 3978 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01875 4540 3993 3980 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01874 3993 3992 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01873 3992 3991 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01872 4540 3990 3992 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01871 3824 3827 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01870 4540 4243 3827 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01869 3697 3832 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01868 3827 3825 3697 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01867 3832 3830 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01866 3830 3828 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01865 4540 3829 3830 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01864 3825 3822 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01863 3822 4261 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01862 4540 4269 3822 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01861 4540 3991 3156 4541 tn L=0.35U W=1.02U AS=0.7854P AD=0.7854P PS=3.6U PD=3.6U 
Mtr_01860 3149 3846 4540 4541 tn L=0.35U W=0.72U AS=0.5544P AD=0.5544P PS=3U PD=3U 
Mtr_01859 3155 3152 3151 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01858 3151 3991 3150 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01857 3150 3156 3154 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01856 3154 3153 3155 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01855 4540 3846 3155 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01854 3148 3149 4540 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01853 3150 3303 3148 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01852 4540 3150 3911 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01851 4540 4243 3305 4541 tn L=0.35U W=1.02U AS=0.7854P AD=0.7854P PS=3.6U PD=3.6U 
Mtr_01850 3304 3983 4540 4541 tn L=0.35U W=0.72U AS=0.5544P AD=0.5544P PS=3U PD=3U 
Mtr_01849 3242 3578 3241 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01848 3241 4243 3308 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01847 3308 3305 3240 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01846 3240 3460 3242 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01845 4540 3983 3242 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01844 3238 3304 4540 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01843 3308 3312 3238 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01842 4540 3308 3303 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01841 4540 3310 3244 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_01840 3244 3327 3316 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_01839 4540 3327 3314 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_01838 3316 3314 3245 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_01837 3245 3313 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_01836 3312 3316 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01835 4540 3578 3313 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01834 3459 4232 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01833 4540 3463 3458 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01832 3461 3458 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01831 3460 3459 3461 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01830 3464 3463 3460 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01829 4540 4232 3464 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01828 3147 3145 3243 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01827 4540 4243 3147 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01826 3143 3144 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01825 3243 3142 3143 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01824 4540 3243 3152 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01823 2865 2868 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01822 4540 4232 2862 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01821 2861 2862 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01820 3145 2865 2861 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01819 2864 4232 3145 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01818 4540 2868 2864 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01817 3237 3239 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01816 4540 4232 3236 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01815 3138 3236 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01814 3142 3237 3138 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01813 3140 4232 3142 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01812 4540 3239 3140 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01811 4540 4107 3037 4541 tn L=0.35U W=1.02U AS=0.7854P AD=0.7854P PS=3.6U PD=3.6U 
Mtr_01810 3039 3035 4540 4541 tn L=0.35U W=0.72U AS=0.5544P AD=0.5544P PS=3U PD=3U 
Mtr_01809 2986 3038 2985 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01808 2985 4107 3042 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01807 3042 3037 2984 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01806 2984 3044 2986 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01805 4540 3035 2986 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01804 2983 3039 4540 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01803 3042 3034 2983 4541 tn L=0.35U W=1.6U AS=1.232P AD=1.232P PS=4.75U PD=4.75U 
Mtr_01802 4540 3042 3153 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01801 4540 2876 2872 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01800 2872 4232 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01799 3034 2869 2872 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01798 2872 4107 3034 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01797 4540 3390 3393 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01796 3391 3390 3295 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01795 3295 3394 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01794 4540 3397 2951 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01793 4540 3390 2965 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01792 2968 3390 2969 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01791 2969 2966 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01790 4540 3397 2964 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01789 2964 3221 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01788 2966 2963 2964 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01787 2964 3226 2966 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01786 4540 3397 2963 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01785 4540 3130 3131 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01784 3130 3390 4540 4541 tn L=0.32U W=0.75U AS=0.5625P AD=0.5625P PS=3U PD=3U 
Mtr_01783 2973 2970 2972 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01782 4540 2973 2974 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01781 2972 2971 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01780 4352 3569 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01779 4540 3570 4352 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01778 4540 3234 3390 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01777 4540 3568 3570 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01776 3401 3404 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01775 3401 3398 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01774 4540 3399 3401 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01773 4540 3401 3397 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01772 4540 3403 3404 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01771 4540 3397 2950 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01770 2950 3380 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01769 2957 2951 2950 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01768 2950 3905 2957 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01767 4540 3390 2956 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01766 2959 3390 2960 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01765 2960 2957 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01764 4540 3397 2954 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01763 4540 3397 2955 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01762 2955 3218 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01761 3127 2954 2955 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01760 2955 3911 3127 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01759 4540 3390 3126 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01758 3128 3390 3024 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01757 3024 3127 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01756 4540 3560 3562 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01755 4540 3567 3561 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01754 4540 3569 3564 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01753 3564 3570 3566 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01752 3566 3561 3565 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01751 3565 3562 3563 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01750 4540 3397 3396 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01749 3296 3396 3394 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01748 3394 3835 3296 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01747 3296 3563 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01746 4540 3651 3557 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01745 3557 3647 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01744 3710 3646 3557 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01743 3557 3799 3710 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01742 3217 3447 3288 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01741 4540 3218 3217 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01740 3216 4458 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01739 3288 3220 3216 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01738 4540 3288 4102 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01737 4198 3382 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01736 4540 3386 3382 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01735 3290 3447 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01734 3382 3380 3290 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01733 3224 3447 3292 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01732 4540 3221 3224 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01731 3223 4470 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01730 3292 3225 3223 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01729 4540 3292 3638 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01728 4540 3641 3544 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01727 3544 3639 3545 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01726 3545 3645 3712 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01725 3640 3643 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_01724 3547 3792 3641 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01723 4540 3640 3547 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01722 4540 3113 3012 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01721 3012 3114 3011 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01720 3011 3112 3991 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01719 4540 3560 3558 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01718 3650 3558 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01717 4540 3559 3650 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01716 3447 3559 4540 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01715 4540 3647 3447 4541 tn L=0.35U W=1.32U AS=1.0164P AD=1.0164P PS=4.2U PD=4.2U 
Mtr_01714 4540 3118 3016 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01713 3016 3389 3015 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01712 3015 3122 3119 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01711 4540 3221 3019 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01710 3019 3553 3120 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01709 4540 3120 3018 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01708 3018 3123 3017 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01707 3017 3119 3635 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01706 3644 3643 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_01705 3551 3907 3642 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01704 4540 3644 3551 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01703 4540 3380 3287 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01702 3287 3553 3379 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01701 4540 3379 3285 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01700 3285 3642 3284 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01699 3284 3378 4196 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01698 4540 4452 3799 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01697 4540 3650 3651 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01696 4540 3646 3220 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01695 4540 3646 3225 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01694 4540 3286 3555 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01693 4540 3559 3554 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01692 4540 3647 3389 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01691 3550 3647 3552 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01690 4540 3550 3553 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01689 3552 3554 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01688 3643 3384 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01687 3384 3383 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01686 4540 3553 3384 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01685 3388 3389 4540 4541 tn L=0.35U W=1.3U AS=1.001P AD=1.001P PS=4.15U PD=4.15U 
Mtr_01684 3294 3445 3646 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01683 4540 3388 3294 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01682 4540 3387 3386 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01681 3291 3445 4540 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01680 3293 3647 3291 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01679 3387 4464 3293 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01678 4540 3289 3215 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01677 3215 3286 3214 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01676 3214 3389 3639 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01675 3114 3115 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01674 3115 3793 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01673 4540 3643 3115 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mtr_01672 4540 3111 3010 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01671 3010 3389 3009 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01670 3009 3117 3112 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01669 3121 3655 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_01668 3020 3555 3122 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01667 4540 3121 3020 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01666 4540 3554 3444 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01665 3444 3555 3445 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01664 3125 3221 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mtr_01663 3023 3553 3124 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01662 4540 3125 3023 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01661 4540 3655 3022 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01660 3022 3555 3021 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01659 3021 3124 3123 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01658 4540 3377 3281 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01657 3281 3376 3280 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01656 3280 3389 3378 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01655 4540 3647 3556 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01654 3556 3650 3645 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01653 4540 3218 3013 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01652 3013 3553 3113 4541 tn L=0.35U W=2.75U AS=2.1175P AD=2.1175P PS=7.05U PD=7.05U 
Mtr_01651 4540 3904 3793 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01650 4540 3793 3014 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mtr_01649 3014 3555 3117 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.n17d 4540 4468 4469 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.n14a 4541 4533 4534 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d0.n18f 4540 4469 4470 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.n16c 4468 4478 4534 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_d0.n15b 4534 4535 4545 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d0.n1 4540 4540 4465 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d0.n14d 4534 4533 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d0.n16d 4534 4478 4468 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_d0.n18d 4540 4469 4470 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.n17a 4469 4468 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.n0 4540 4540 4466 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d0.n4b 4540 4467 4494 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d0.n16a 4468 4478 4534 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_d0.n16b 4534 4478 4468 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_d0.n15c 4545 4535 4534 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d0.n17b 4540 4468 4469 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.n18a 4470 4469 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.n6d 4532 4494 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d0.n3 4465 4466 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d0.n7d 4541 4493 4533 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d0.n5a 4493 4465 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d0.n7c 4533 4493 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d0.n18e 4470 4469 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.n6c 4541 4494 4532 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d0.n14b 4534 4533 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d0.n6b 4532 4494 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d0.n7b 4541 4493 4533 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d0.n15a 4545 4535 4534 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d0.n7a 4533 4493 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d0.n6a 4541 4494 4532 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d0.n8d 4532 4535 4531 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d0.n8c 4531 4535 4532 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d0.n8b 4532 4535 4531 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d0.n8a 4531 4535 4532 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d0.n18b 4540 4469 4470 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.n4a 4494 4467 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d0.n17c 4469 4468 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d0.n14c 4541 4533 4534 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d0.n15d 4534 4535 4545 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d0.n2 4465 4540 4467 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d0.n5b 4540 4465 4493 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d0.n18c 4470 4469 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.n17d 4540 4462 4463 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.n14a 4541 4528 4529 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d1.n18f 4540 4463 4464 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.n16c 4462 4478 4529 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_d1.n15b 4529 4535 4544 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d1.n1 4540 4540 4459 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d1.n14d 4529 4528 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d1.n16d 4529 4478 4462 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_d1.n18d 4540 4463 4464 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.n17a 4463 4462 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.n0 4540 4540 4460 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d1.n4b 4540 4461 4492 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d1.n16a 4462 4478 4529 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_d1.n16b 4529 4478 4462 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_d1.n15c 4544 4535 4529 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d1.n17b 4540 4462 4463 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.n18a 4464 4463 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.n6d 4526 4492 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d1.n3 4459 4460 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d1.n7d 4541 4491 4528 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d1.n5a 4491 4459 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d1.n7c 4528 4491 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d1.n18e 4464 4463 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.n6c 4541 4492 4526 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d1.n14b 4529 4528 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d1.n6b 4526 4492 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d1.n7b 4541 4491 4528 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d1.n15a 4544 4535 4529 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d1.n7a 4528 4491 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d1.n6a 4541 4492 4526 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d1.n8d 4526 4535 4527 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d1.n8c 4527 4535 4526 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d1.n8b 4526 4535 4527 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d1.n8a 4527 4535 4526 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d1.n18b 4540 4463 4464 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.n4a 4492 4461 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d1.n17c 4463 4462 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d1.n14c 4541 4528 4529 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d1.n15d 4529 4535 4544 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d1.n2 4459 4540 4461 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d1.n5b 4540 4459 4491 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d1.n18c 4464 4463 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.n17d 4540 60 61 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.n14a 4541 10 59 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i7.n18f 4540 61 123 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.n16c 60 4478 59 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i7.n15b 59 4535 9 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i7.n1 4540 4540 57 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i7.n14d 59 10 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i7.n16d 59 4478 60 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i7.n18d 4540 61 123 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.n17a 61 60 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.n0 4540 4540 55 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i7.n4b 4540 56 58 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i7.n16a 60 4478 59 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i7.n16b 59 4478 60 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i7.n15c 9 4535 59 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i7.n17b 4540 60 61 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.n18a 123 61 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.n6d 8 58 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i7.n3 57 55 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i7.n7d 4541 54 10 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i7.n5a 54 57 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i7.n7c 10 54 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i7.n18e 123 61 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.n6c 4541 58 8 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i7.n14b 59 10 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i7.n6b 8 58 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i7.n7b 4541 54 10 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i7.n15a 9 4535 59 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i7.n7a 10 54 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i7.n6a 4541 58 8 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i7.n8d 8 4535 6 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i7.n8c 6 4535 8 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i7.n8b 8 4535 6 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i7.n8a 6 4535 8 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i7.n18b 4540 61 123 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.n4a 58 56 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i7.n17c 61 60 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i7.n14c 4541 10 59 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i7.n15d 59 4535 9 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i7.n2 57 4540 56 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i7.n5b 4540 57 54 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i7.n18c 123 61 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.n16b 4540 4478 1663 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_ovr.n1 4540 3715 1830 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_ovr.n17a 1662 1663 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.n18d 4540 1662 1550 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.n14d 1549 1694 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ovr.n16d 4540 4478 1663 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_ovr.n16a 1663 4478 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_ovr.n15b 1549 4535 1828 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ovr.n14a 4541 1694 1549 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ovr.n16c 1663 4478 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_ovr.n18f 4540 1662 1550 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.n18c 1550 1662 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.n17d 4540 1663 1662 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.n5b 4540 1830 1832 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_ovr.n14c 4541 1694 1549 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ovr.n2 1830 4478 1829 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_ovr.n15d 1549 4535 1828 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ovr.n18b 4540 1662 1550 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.n17c 1662 1663 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.n8a 1942 4535 1693 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ovr.n8b 1693 4535 1942 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ovr.n8c 1942 4535 1693 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ovr.n8d 1693 4535 1942 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ovr.n6a 4541 1695 1693 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ovr.n14b 1549 1694 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ovr.n7a 1694 1832 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ovr.n15a 1828 4535 1549 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ovr.n4a 1695 1829 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_ovr.n5a 1832 1830 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_ovr.n7b 4541 1832 1694 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ovr.n3 1830 1831 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_ovr.n6b 1693 1695 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ovr.n6c 4541 1695 1693 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ovr.n18a 1550 1662 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.n7c 1694 1832 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ovr.n18e 1550 1662 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.n7d 4541 1832 1694 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ovr.n17b 4540 1663 1662 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ovr.n6d 1693 1695 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ovr.n15c 1828 4535 1549 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ovr.n4b 4540 1829 1695 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_ovr.n0 4540 4478 1831 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y0.n18c 4443 4442 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.n14a 4541 4513 4514 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y0.n15b 4514 4535 4539 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y0.n16c 4441 4478 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_y0.n1 4540 4436 4438 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y0.n14d 4514 4513 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y0.n18d 4540 4442 4443 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.n16d 4540 4478 4441 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_y0.n17a 4442 4441 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.n16a 4441 4478 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_y0.n4b 4540 4440 4486 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y0.n0 4540 4437 4439 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y0.n16b 4540 4478 4441 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_y0.n6d 4512 4486 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y0.n15c 4539 4535 4514 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y0.n7d 4541 4485 4513 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y0.n17b 4540 4441 4442 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.n7c 4513 4485 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y0.n4a 4486 4440 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y0.n6c 4541 4486 4512 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y0.n6b 4512 4486 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y0.n18e 4443 4442 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.n18a 4443 4442 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.n3 4438 4439 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y0.n7b 4541 4485 4513 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y0.n7a 4513 4485 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y0.n5a 4485 4438 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y0.n6a 4541 4486 4512 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y0.n15a 4539 4535 4514 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y0.n8d 4512 4535 4511 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y0.n14b 4514 4513 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y0.n8c 4511 4535 4512 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y0.n8b 4512 4535 4511 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y0.n8a 4511 4535 4512 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y0.n17c 4442 4441 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.n2 4438 4437 4440 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y0.n18b 4540 4442 4443 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.n15d 4514 4535 4539 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y0.n18f 4540 4442 4443 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y0.n14c 4541 4513 4514 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y0.n5b 4540 4438 4485 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y0.n17d 4540 4441 4442 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.n17d 4540 1278 1398 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.n14a 4541 1400 1401 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b0.n18f 4540 1398 1399 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.n16c 1278 4478 1401 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_b0.n15b 1401 4535 1402 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b0.n1 4540 4540 993 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b0.n14d 1401 1400 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b0.n16d 1401 4478 1278 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_b0.n18d 4540 1398 1399 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.n17a 1398 1278 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.n0 4540 4540 994 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b0.n4b 4540 1104 1240 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b0.n16a 1278 4478 1401 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_b0.n16b 1401 4478 1278 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_b0.n15c 1402 4535 1401 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b0.n17b 4540 1278 1398 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.n18a 1399 1398 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.n6d 1241 1240 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b0.n3 993 994 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b0.n7d 4541 1239 1400 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b0.n5a 1239 993 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b0.n7c 1400 1239 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b0.n18e 1399 1398 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.n6c 4541 1240 1241 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b0.n14b 1401 1400 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b0.n6b 1241 1240 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b0.n7b 4541 1239 1400 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b0.n15a 1402 4535 1401 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b0.n7a 1400 1239 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b0.n6a 4541 1240 1241 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b0.n8d 1241 4535 1242 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b0.n8c 1242 4535 1241 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b0.n8b 1241 4535 1242 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b0.n8a 1242 4535 1241 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b0.n18b 4540 1398 1399 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.n4a 1240 1104 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b0.n17c 1398 1278 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b0.n14c 4541 1400 1401 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b0.n15d 1401 4535 1402 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b0.n2 993 4540 1104 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b0.n5b 4540 993 1239 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b0.n18c 1399 1398 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.n17d 4540 3572 3660 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.n14a 4541 3686 3687 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a0.n18f 4540 3660 3661 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.n16c 3572 4478 3687 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_a0.n15b 3687 4535 3662 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a0.n1 4540 4540 3405 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a0.n14d 3687 3686 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a0.n16d 3687 4478 3572 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_a0.n18d 4540 3660 3661 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.n17a 3660 3572 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.n0 4540 4540 3300 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a0.n4b 4540 3406 3451 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a0.n16a 3572 4478 3687 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_a0.n16b 3687 4478 3572 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_a0.n15c 3662 4535 3687 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a0.n17b 4540 3572 3660 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.n18a 3661 3660 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.n6d 3454 3451 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a0.n3 3405 3300 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a0.n7d 4541 3450 3686 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a0.n5a 3450 3405 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a0.n7c 3686 3450 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a0.n18e 3661 3660 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.n6c 4541 3451 3454 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a0.n14b 3687 3686 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a0.n6b 3454 3451 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a0.n7b 4541 3450 3686 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a0.n15a 3662 4535 3687 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a0.n7a 3686 3450 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a0.n6a 4541 3451 3454 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a0.n8d 3454 4535 3453 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a0.n8c 3453 4535 3454 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a0.n8b 3454 4535 3453 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a0.n8a 3453 4535 3454 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a0.n18b 4540 3660 3661 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.n4a 3451 3406 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a0.n17c 3660 3572 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a0.n14c 4541 3686 3687 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a0.n15d 3687 4535 3662 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a0.n2 3405 4540 3406 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a0.n5b 4540 3405 3450 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a0.n18c 3661 3660 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vsseck1.75onymous_ 4540 4473 4445 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vsseck1.39onymous_ 4540 4476 4474 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vsseck1.13onymous_ 4540 4474 4445 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vsseck1.34onymous_ 4445 4474 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vsseck1.65onymous_ 4445 4473 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vsseck1.91onymous_ 4473 4476 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vsseck1.28onymous_ 4540 4474 4445 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vsseck1.86onymous_ 4540 4473 4445 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vsseck1.23onymous_ 4445 4474 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vsseck1.80onymous_ 4445 4473 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.n14c 4541 4366 4358 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_r3.n6d 4365 4364 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r3.n15d 4358 4535 4371 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_r3.n5b 4540 4373 4374 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_r3.n18c 4350 4355 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.n17d 4540 4359 4355 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.n14a 4541 4366 4358 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_r3.n16c 4359 4478 4358 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_r3.n18f 4540 4355 4350 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.n15b 4358 4535 4371 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_r3.n1 4540 4368 4373 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_r3.n16d 4358 4478 4359 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_r3.n14d 4358 4366 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_r3.n18d 4540 4355 4350 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.n17a 4355 4359 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.n4b 4540 4367 4364 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_r3.n0 4540 4372 4375 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_r3.n16a 4359 4478 4358 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_r3.n4a 4364 4367 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_r3.n16b 4358 4478 4359 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_r3.n15c 4371 4535 4358 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_r3.n17b 4540 4359 4355 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.n18a 4350 4355 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.n3 4373 4375 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_r3.n7d 4541 4374 4366 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r3.n5a 4374 4373 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_r3.n7c 4366 4374 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r3.n18e 4350 4355 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.n6c 4541 4364 4365 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r3.n14b 4358 4366 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_r3.n6b 4365 4364 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r3.n7b 4541 4374 4366 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r3.n15a 4371 4535 4358 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_r3.n7a 4366 4374 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r3.n6a 4541 4364 4365 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r3.n8d 4365 4535 4370 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r3.n8c 4370 4535 4365 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r3.n8b 4365 4535 4370 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r3.n8a 4370 4535 4365 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r3.n2 4373 4372 4367 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_r3.n18b 4540 4355 4350 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r3.n17c 4355 4359 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.n14c 4541 4081 3971 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_q3.n6d 4080 4079 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q3.n15d 3971 4535 4128 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_q3.n5b 4540 4129 4130 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_q3.n18c 4071 3933 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.n17d 4540 3970 3933 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.n14a 4541 4081 3971 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_q3.n16c 3970 4478 3971 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_q3.n18f 4540 3933 4071 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.n15b 3971 4535 4128 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_q3.n1 4540 4084 4129 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_q3.n16d 3971 4478 3970 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_q3.n14d 3971 4081 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_q3.n18d 4540 3933 4071 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.n17a 3933 3970 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.n4b 4540 4082 4079 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_q3.n0 4540 4121 4083 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_q3.n16a 3970 4478 3971 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_q3.n4a 4079 4082 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_q3.n16b 3971 4478 3970 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_q3.n15c 4128 4535 3971 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_q3.n17b 4540 3970 3933 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.n18a 4071 3933 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.n3 4129 4083 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_q3.n7d 4541 4130 4081 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q3.n5a 4130 4129 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_q3.n7c 4081 4130 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q3.n18e 4071 3933 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.n6c 4541 4079 4080 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q3.n14b 3971 4081 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_q3.n6b 4080 4079 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q3.n7b 4541 4130 4081 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q3.n15a 4128 4535 3971 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_q3.n7a 4081 4130 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q3.n6a 4541 4079 4080 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q3.n8d 4080 4535 4126 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q3.n8c 4126 4535 4080 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q3.n8b 4080 4535 4126 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q3.n8a 4126 4535 4080 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q3.n2 4129 4121 4082 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_q3.n18b 4540 3933 4071 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q3.n17c 3933 3970 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.n18c 4419 4418 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.n14a 4541 4498 4499 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y3.n15b 4499 4535 4536 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y3.n16c 4417 4478 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_y3.n1 4540 4412 4414 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y3.n14d 4499 4498 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y3.n18d 4540 4418 4419 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.n16d 4540 4478 4417 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_y3.n17a 4418 4417 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.n16a 4417 4478 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_y3.n4b 4540 4416 4480 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y3.n0 4540 4413 4415 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y3.n16b 4540 4478 4417 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_y3.n6d 4497 4480 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y3.n15c 4536 4535 4499 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y3.n7d 4541 4479 4498 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y3.n17b 4540 4417 4418 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.n7c 4498 4479 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y3.n4a 4480 4416 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y3.n6c 4541 4480 4497 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y3.n6b 4497 4480 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y3.n18e 4419 4418 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.n18a 4419 4418 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.n3 4414 4415 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y3.n7b 4541 4479 4498 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y3.n7a 4498 4479 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y3.n5a 4479 4414 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y3.n6a 4541 4480 4497 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y3.n15a 4536 4535 4499 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y3.n8d 4497 4535 4496 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y3.n14b 4499 4498 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y3.n8c 4496 4535 4497 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y3.n8b 4497 4535 4496 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y3.n8a 4496 4535 4497 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y3.n17c 4418 4417 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.n2 4414 4413 4416 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y3.n18b 4540 4418 4419 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.n15d 4499 4535 4536 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y3.n18f 4540 4418 4419 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y3.n14c 4541 4498 4499 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y3.n5b 4540 4414 4479 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y3.n17d 4540 4417 4418 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.n16b 4540 4478 2860 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_np.n1 4540 3188 3028 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_np.n17a 2754 2860 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.n18d 4540 2754 2717 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.n14d 2753 2981 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_np.n16d 4540 4478 2860 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_np.n16a 2860 4478 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_np.n15b 2753 4535 3027 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_np.n14a 4541 2981 2753 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_np.n16c 2860 4478 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_np.n18f 4540 2754 2717 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.n18c 2717 2754 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.n17d 4540 2860 2754 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.n5b 4540 3028 3030 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_np.n14c 4541 2981 2753 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_np.n2 3028 4478 2982 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_np.n15d 2753 4535 3027 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_np.n18b 4540 2754 2717 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.n17c 2754 2860 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.n8a 3026 4535 2980 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_np.n8b 2980 4535 3026 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_np.n8c 3026 4535 2980 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_np.n8d 2980 4535 3026 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_np.n6a 4541 2979 2980 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_np.n14b 2753 2981 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_np.n7a 2981 3030 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_np.n15a 3027 4535 2753 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_np.n4a 2979 2982 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_np.n5a 3030 3028 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_np.n7b 4541 3030 2981 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_np.n3 3028 3029 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_np.n6b 2980 2979 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_np.n6c 4541 2979 2980 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_np.n18a 2717 2754 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.n7c 2981 3030 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_np.n18e 2717 2754 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.n7d 4541 3030 2981 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_np.n17b 4540 2860 2754 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_np.n6d 2980 2979 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_np.n15c 3027 4535 2753 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_np.n4b 4540 2982 2979 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_np.n0 4540 4478 3029 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_ck.n18a 4476 172 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ck.n16b 173 4478 174 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_ck.n17c 172 174 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ck.n18f 4540 172 4476 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ck.n14b 173 169 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ck.n14c 4541 169 173 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ck.n17a 172 174 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ck.n18e 4476 172 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ck.n15c 180 4535 173 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ck.n17d 4540 174 172 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ck.n18b 4540 172 4476 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ck.n14d 173 169 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ck.n6d 168 4541 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ck.n7d 4541 4535 169 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ck.n7c 169 4535 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ck.n6c 4541 4541 168 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ck.n16c 174 4478 173 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_ck.n6b 168 4541 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ck.n7b 4541 4535 169 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ck.n7a 169 4535 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ck.n6a 4541 4541 168 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ck.n15a 180 4535 173 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ck.n8d 168 4535 178 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ck.n8c 178 4535 168 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ck.n18c 4476 172 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ck.n8b 168 4535 178 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ck.n16d 173 4478 174 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_ck.n8a 178 4535 168 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ck.n15d 173 4535 180 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ck.n14a 4541 169 173 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ck.n18d 4540 172 4476 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ck.n16a 174 4478 173 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_ck.n17b 4540 174 172 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ck.n15b 173 4535 180 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i2.n17d 4540 104 105 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.n14a 4541 35 103 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i2.n18f 4540 105 3647 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.n16c 104 4478 103 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i2.n15b 103 4535 34 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i2.n1 4540 4540 100 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i2.n14d 103 35 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i2.n16d 103 4478 104 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i2.n18d 4540 105 3647 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.n17a 105 104 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.n0 4540 4540 99 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i2.n4b 4540 101 102 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i2.n16a 104 4478 103 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i2.n16b 103 4478 104 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i2.n15c 34 4535 103 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i2.n17b 4540 104 105 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.n18a 3647 105 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.n6d 33 102 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i2.n3 100 99 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i2.n7d 4541 98 35 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i2.n5a 98 100 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i2.n7c 35 98 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i2.n18e 3647 105 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.n6c 4541 102 33 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i2.n14b 103 35 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i2.n6b 33 102 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i2.n7b 4541 98 35 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i2.n15a 34 4535 103 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i2.n7a 35 98 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i2.n6a 4541 102 33 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i2.n8d 33 4535 31 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i2.n8c 31 4535 33 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i2.n8b 33 4535 31 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i2.n8a 31 4535 33 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i2.n18b 4540 105 3647 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.n4a 102 101 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i2.n17c 105 104 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i2.n14c 4541 35 103 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i2.n15d 103 4535 34 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i2.n2 100 4540 101 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i2.n5b 4540 100 98 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i2.n18c 3647 105 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.n16b 4540 4478 139 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_f3.n1 4540 148 152 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_f3.n17a 136 139 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.n18d 4540 136 132 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.n14d 135 146 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_f3.n16d 4540 4478 139 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_f3.n16a 139 4478 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_f3.n15b 135 4535 151 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_f3.n14a 4541 146 135 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_f3.n16c 139 4478 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_f3.n18f 4540 136 132 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.n18c 132 136 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.n17d 4540 139 136 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.n5b 4540 152 154 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_f3.n14c 4541 146 135 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_f3.n2 152 4478 147 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_f3.n15d 135 4535 151 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_f3.n18b 4540 136 132 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.n17c 136 139 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.n8a 150 4535 145 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_f3.n8b 145 4535 150 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_f3.n8c 150 4535 145 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_f3.n8d 145 4535 150 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_f3.n6a 4541 144 145 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_f3.n14b 135 146 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_f3.n7a 146 154 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_f3.n15a 151 4535 135 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_f3.n4a 144 147 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_f3.n5a 154 152 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_f3.n7b 4541 154 146 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_f3.n3 152 153 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_f3.n6b 145 144 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_f3.n6c 4541 144 145 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_f3.n18a 132 136 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.n7c 146 154 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_f3.n18e 132 136 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.n7d 4541 154 146 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_f3.n17b 4540 139 136 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_f3.n6d 145 144 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_f3.n15c 151 4535 135 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_f3.n4b 4540 147 144 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_f3.n0 4540 4478 153 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_zero.n16b 4540 4478 1106 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_zero.n1 4540 2790 1281 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_zero.n17a 996 1106 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.n18d 4540 996 952 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.n14d 995 1245 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_zero.n16d 4540 4478 1106 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_zero.n16a 1106 4478 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_zero.n15b 995 4535 1280 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_zero.n14a 4541 1245 995 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_zero.n16c 1106 4478 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_zero.n18f 4540 996 952 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.n18c 952 996 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.n17d 4540 1106 996 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.n5b 4540 1281 1283 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_zero.n14c 4541 1245 995 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_zero.n2 1281 4478 1246 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_zero.n15d 995 4535 1280 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_zero.n18b 4540 996 952 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.n17c 996 1106 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.n8a 1279 4535 1244 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_zero.n8b 1244 4535 1279 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_zero.n8c 1279 4535 1244 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_zero.n8d 1244 4535 1279 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_zero.n6a 4541 1243 1244 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_zero.n14b 995 1245 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_zero.n7a 1245 1283 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_zero.n15a 1280 4535 995 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_zero.n4a 1243 1246 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_zero.n5a 1283 1281 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_zero.n7b 4541 1283 1245 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_zero.n3 1281 1282 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_zero.n6b 1244 1243 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_zero.n6c 4541 1243 1244 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_zero.n18a 952 996 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.n7c 1245 1283 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_zero.n18e 952 996 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.n7d 4541 1283 1245 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_zero.n17b 4540 1106 996 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_zero.n6d 1244 1243 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_zero.n15c 1280 4535 995 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_zero.n4b 4540 1246 1243 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_zero.n0 4540 4478 1282 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i3.n17d 4540 96 97 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.n14a 4541 30 95 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i3.n18f 4540 97 130 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.n16c 96 4478 95 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i3.n15b 95 4535 29 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i3.n1 4540 4540 94 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i3.n14d 95 30 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i3.n16d 95 4478 96 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i3.n18d 4540 97 130 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.n17a 97 96 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.n0 4540 4540 91 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i3.n4b 4540 93 92 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i3.n16a 96 4478 95 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i3.n16b 95 4478 96 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i3.n15c 29 4535 95 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i3.n17b 4540 96 97 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.n18a 130 97 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.n6d 28 92 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i3.n3 94 91 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i3.n7d 4541 90 30 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i3.n5a 90 94 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i3.n7c 30 90 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i3.n18e 130 97 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.n6c 4541 92 28 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i3.n14b 95 30 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i3.n6b 28 92 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i3.n7b 4541 90 30 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i3.n15a 29 4535 95 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i3.n7a 30 90 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i3.n6a 4541 92 28 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i3.n8d 28 4535 26 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i3.n8c 26 4535 28 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i3.n8b 28 4535 26 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i3.n8a 26 4535 28 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i3.n18b 4540 97 130 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.n4a 92 93 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i3.n17c 97 96 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i3.n14c 4541 30 95 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i3.n15d 95 4535 29 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i3.n2 94 4540 93 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i3.n5b 4540 94 90 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i3.n18c 130 97 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddeck1.38onymous_ 4540 79 126 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddeck1.64onymous_ 4540 4476 79 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddeck1.116nymous_ 78 4476 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddeck1.90onymous_ 126 78 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddeck1.59onymous_ 126 79 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddeck1.111nymous_ 4540 78 126 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddeck1.53onymous_ 4540 79 126 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddeck1.48onymous_ 126 79 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddeck1.105nymous_ 126 78 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddeck1.100nymous_ 4540 78 126 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.n14c 4541 4378 4379 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_r0.n6d 4363 4361 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r0.n15d 4379 4535 4380 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_r0.n5b 4540 4354 4360 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_r0.n18c 4377 4376 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.n17d 4540 4369 4376 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.n14a 4541 4378 4379 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_r0.n16c 4369 4478 4379 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_r0.n18f 4540 4376 4377 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.n15b 4379 4535 4380 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_r0.n1 4540 4351 4354 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_r0.n16d 4379 4478 4369 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_r0.n14d 4379 4378 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_r0.n18d 4540 4376 4377 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.n17a 4376 4369 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.n4b 4540 4356 4361 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_r0.n0 4540 4352 4353 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_r0.n16a 4369 4478 4379 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_r0.n4a 4361 4356 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_r0.n16b 4379 4478 4369 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_r0.n15c 4380 4535 4379 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_r0.n17b 4540 4369 4376 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.n18a 4377 4376 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.n3 4354 4353 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_r0.n7d 4541 4360 4378 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r0.n5a 4360 4354 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_r0.n7c 4378 4360 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r0.n18e 4377 4376 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.n6c 4541 4361 4363 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r0.n14b 4379 4378 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_r0.n6b 4363 4361 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r0.n7b 4541 4360 4378 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r0.n15a 4380 4535 4379 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_r0.n7a 4378 4360 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r0.n6a 4541 4361 4363 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r0.n8d 4363 4535 4362 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r0.n8c 4362 4535 4363 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r0.n8b 4363 4535 4362 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r0.n8a 4362 4535 4363 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_r0.n2 4354 4352 4356 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_r0.n18b 4540 4376 4377 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_r0.n17c 4376 4369 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.n14c 4541 4230 4231 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_q0.n6d 4078 4075 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q0.n15d 4231 4535 4125 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_q0.n5b 4540 3932 4076 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_q0.n18c 4342 4229 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.n17d 4540 4124 4229 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.n14a 4541 4230 4231 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_q0.n16c 4124 4478 4231 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_q0.n18f 4540 4229 4342 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.n15b 4231 4535 4125 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_q0.n1 4540 3931 3932 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_q0.n16d 4231 4478 4124 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_q0.n14d 4231 4230 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_q0.n18d 4540 4229 4342 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.n17a 4229 4124 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.n4b 4540 3968 4075 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_q0.n0 4540 4352 3930 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_q0.n16a 4124 4478 4231 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_q0.n4a 4075 3968 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_q0.n16b 4231 4478 4124 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_q0.n15c 4125 4535 4231 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_q0.n17b 4540 4124 4229 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.n18a 4342 4229 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.n3 3932 3930 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_q0.n7d 4541 4076 4230 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q0.n5a 4076 3932 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_q0.n7c 4230 4076 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q0.n18e 4342 4229 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.n6c 4541 4075 4078 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q0.n14b 4231 4230 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_q0.n6b 4078 4075 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q0.n7b 4541 4076 4230 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q0.n15a 4125 4535 4231 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_q0.n7a 4230 4076 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q0.n6a 4541 4075 4078 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q0.n8d 4078 4535 4077 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q0.n8c 4077 4535 4078 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q0.n8b 4078 4535 4077 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q0.n8a 4077 4535 4078 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_q0.n2 3932 4352 3968 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_q0.n18b 4540 4229 4342 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_q0.n17c 4229 4124 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vssick0.31onymous_ 4444 4471 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vssick0.25onymous_ 4540 4471 4444 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vssick0.81onymous_ 4540 4472 4444 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vssick0.75onymous_ 4444 4472 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vssick0.46onymous_ 4444 4471 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vssick0.20onymous_ 4471 4476 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vssick0.70onymous_ 4540 4476 4472 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vssick0.96onymous_ 4540 4472 4444 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vssick0.36onymous_ 4540 4471 4444 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vssick0.86onymous_ 4444 4472 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.n17d 4540 149 155 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.n14a 4541 157 158 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b3.n18f 4540 155 156 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.n16c 149 4478 158 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_b3.n15b 158 4535 159 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b3.n1 4540 4540 133 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b3.n14d 158 157 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b3.n16d 158 4478 149 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_b3.n18d 4540 155 156 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.n17a 155 149 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.n0 4540 4540 134 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b3.n4b 4540 137 141 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b3.n16a 149 4478 158 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_b3.n16b 158 4478 149 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_b3.n15c 159 4535 158 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b3.n17b 4540 149 155 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.n18a 156 155 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.n6d 142 141 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b3.n3 133 134 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b3.n7d 4541 140 157 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b3.n5a 140 133 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b3.n7c 157 140 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b3.n18e 156 155 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.n6c 4541 141 142 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b3.n14b 158 157 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b3.n6b 142 141 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b3.n7b 4541 140 157 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b3.n15a 159 4535 158 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b3.n7a 157 140 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b3.n6a 4541 141 142 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b3.n8d 142 4535 143 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b3.n8c 143 4535 142 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b3.n8b 142 4535 143 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b3.n8a 143 4535 142 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b3.n18b 4540 155 156 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.n4a 141 137 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b3.n17c 155 149 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b3.n14c 4541 157 158 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b3.n15d 158 4535 159 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b3.n2 133 4540 137 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b3.n5b 4540 133 140 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b3.n18c 156 155 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.n17d 4540 1826 1940 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.n14a 4541 1970 1971 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a3.n18f 4540 1940 2930 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.n16c 1826 4478 1971 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_a3.n15b 1971 4535 1941 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a3.n1 4540 4540 1660 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a3.n14d 1971 1970 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a3.n16d 1971 4478 1826 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_a3.n18d 4540 1940 2930 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.n17a 1940 1826 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.n0 4540 4540 1548 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a3.n4b 4540 1661 1689 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a3.n16a 1826 4478 1971 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_a3.n16b 1971 4478 1826 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_a3.n15c 1941 4535 1971 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a3.n17b 4540 1826 1940 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.n18a 2930 1940 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.n6d 1692 1689 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a3.n3 1660 1548 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a3.n7d 4541 1827 1970 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a3.n5a 1827 1660 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a3.n7c 1970 1827 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a3.n18e 2930 1940 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.n6c 4541 1689 1692 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a3.n14b 1971 1970 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a3.n6b 1692 1689 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a3.n7b 4541 1827 1970 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a3.n15a 1941 4535 1971 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a3.n7a 1970 1827 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a3.n6a 4541 1689 1692 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a3.n8d 1692 4535 1691 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a3.n8c 1691 4535 1692 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a3.n8b 1692 4535 1691 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a3.n8a 1691 4535 1692 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a3.n18b 4540 1940 2930 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.n4a 1689 1661 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a3.n17c 1940 1826 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a3.n14c 4541 1970 1971 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a3.n15d 1971 4535 1941 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a3.n2 1660 4540 1661 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a3.n5b 4540 1660 1827 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a3.n18c 2930 1940 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.n17d 4540 4456 4457 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.n14a 4541 4523 4524 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d2.n18f 4540 4457 4458 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.n16c 4456 4478 4524 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_d2.n15b 4524 4535 4543 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d2.n1 4540 4540 4454 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d2.n14d 4524 4523 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d2.n16d 4524 4478 4456 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_d2.n18d 4540 4457 4458 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.n17a 4457 4456 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.n0 4540 4540 4453 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d2.n4b 4540 4455 4489 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d2.n16a 4456 4478 4524 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_d2.n16b 4524 4478 4456 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_d2.n15c 4543 4535 4524 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d2.n17b 4540 4456 4457 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.n18a 4458 4457 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.n6d 4522 4489 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d2.n3 4454 4453 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d2.n7d 4541 4490 4523 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d2.n5a 4490 4454 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d2.n7c 4523 4490 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d2.n18e 4458 4457 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.n6c 4541 4489 4522 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d2.n14b 4524 4523 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d2.n6b 4522 4489 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d2.n7b 4541 4490 4523 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d2.n15a 4543 4535 4524 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d2.n7a 4523 4490 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d2.n6a 4541 4489 4522 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d2.n8d 4522 4535 4521 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d2.n8c 4521 4535 4522 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d2.n8b 4522 4535 4521 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d2.n8a 4521 4535 4522 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d2.n18b 4540 4457 4458 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.n4a 4489 4455 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d2.n17c 4457 4456 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d2.n14c 4541 4523 4524 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d2.n15d 4524 4535 4543 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d2.n2 4454 4540 4455 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d2.n5b 4540 4454 4490 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d2.n18c 4458 4457 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.n17d 4540 52 53 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.n14a 4541 5 51 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i8.n18f 4540 53 122 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.n16c 52 4478 51 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i8.n15b 51 4535 4 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i8.n1 4540 4540 47 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i8.n14d 51 5 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i8.n16d 51 4478 52 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i8.n18d 4540 53 122 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.n17a 53 52 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.n0 4540 4540 48 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i8.n4b 4540 49 50 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i8.n16a 52 4478 51 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i8.n16b 51 4478 52 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i8.n15c 4 4535 51 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i8.n17b 4540 52 53 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.n18a 122 53 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.n6d 3 50 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i8.n3 47 48 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i8.n7d 4541 46 5 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i8.n5a 46 47 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i8.n7c 5 46 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i8.n18e 122 53 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.n6c 4541 50 3 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i8.n14b 51 5 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i8.n6b 3 50 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i8.n7b 4541 46 5 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i8.n15a 4 4535 51 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i8.n7a 5 46 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i8.n6a 4541 50 3 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i8.n8d 3 4535 1 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i8.n8c 1 4535 3 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i8.n8b 3 4535 1 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i8.n8a 1 4535 3 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i8.n18b 4540 53 122 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.n4a 50 49 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i8.n17c 53 52 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i8.n14c 4541 5 51 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i8.n15d 51 4535 4 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i8.n2 47 4540 49 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i8.n5b 4540 47 46 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i8.n18c 122 53 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.n18c 4435 4434 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.n14a 4541 4508 4509 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y1.n15b 4509 4535 4538 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y1.n16c 4433 4478 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_y1.n1 4540 4429 4431 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y1.n14d 4509 4508 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y1.n18d 4540 4434 4435 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.n16d 4540 4478 4433 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_y1.n17a 4434 4433 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.n16a 4433 4478 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_y1.n4b 4540 4432 4483 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y1.n0 4540 4430 4428 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y1.n16b 4540 4478 4433 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_y1.n6d 4506 4483 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y1.n15c 4538 4535 4509 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y1.n7d 4541 4484 4508 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y1.n17b 4540 4433 4434 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.n7c 4508 4484 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y1.n4a 4483 4432 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y1.n6c 4541 4483 4506 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y1.n6b 4506 4483 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y1.n18e 4435 4434 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.n18a 4435 4434 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.n3 4431 4428 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y1.n7b 4541 4484 4508 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y1.n7a 4508 4484 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y1.n5a 4484 4431 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y1.n6a 4541 4483 4506 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y1.n15a 4538 4535 4509 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y1.n8d 4506 4535 4507 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y1.n14b 4509 4508 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y1.n8c 4507 4535 4506 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y1.n8b 4506 4535 4507 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y1.n8a 4507 4535 4506 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y1.n17c 4434 4433 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.n2 4431 4430 4432 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y1.n18b 4540 4434 4435 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.n15d 4509 4535 4538 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y1.n18f 4540 4434 4435 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y1.n14c 4541 4508 4509 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y1.n5b 4540 4431 4484 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y1.n17d 4540 4433 4434 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddeck0.38onymous_ 4540 81 127 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddeck0.64onymous_ 4540 4476 81 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddeck0.116nymous_ 80 4476 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddeck0.90onymous_ 127 80 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddeck0.59onymous_ 127 81 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddeck0.111nymous_ 4540 80 127 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddeck0.53onymous_ 4540 81 127 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddeck0.48onymous_ 127 81 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddeck0.105nymous_ 127 80 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddeck0.100nymous_ 4540 80 127 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.n17d 4540 88 89 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.n14a 4541 25 87 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i4.n18f 4540 89 128 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.n16c 88 4478 87 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i4.n15b 87 4535 24 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i4.n1 4540 4540 83 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i4.n14d 87 25 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i4.n16d 87 4478 88 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i4.n18d 4540 89 128 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.n17a 89 88 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.n0 4540 4540 84 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i4.n4b 4540 85 86 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i4.n16a 88 4478 87 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i4.n16b 87 4478 88 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i4.n15c 24 4535 87 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i4.n17b 4540 88 89 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.n18a 128 89 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.n6d 23 86 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i4.n3 83 84 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i4.n7d 4541 82 25 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i4.n5a 82 83 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i4.n7c 25 82 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i4.n18e 128 89 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.n6c 4541 86 23 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i4.n14b 87 25 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i4.n6b 23 86 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i4.n7b 4541 82 25 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i4.n15a 24 4535 87 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i4.n7a 25 82 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i4.n6a 4541 86 23 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i4.n8d 23 4535 21 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i4.n8c 21 4535 23 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i4.n8b 23 4535 21 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i4.n8a 21 4535 23 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i4.n18b 4540 89 128 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.n4a 86 85 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i4.n17c 89 88 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i4.n14c 4541 25 87 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i4.n15d 87 4535 24 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i4.n2 83 4540 85 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i4.n5b 4540 83 82 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i4.n18c 128 89 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.n17d 4540 170 175 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.n14a 4541 200 201 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b2.n18f 4540 175 176 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.n16c 170 4478 201 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_b2.n15b 201 4535 177 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b2.n1 4540 4540 162 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b2.n14d 201 200 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b2.n16d 201 4478 170 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_b2.n18d 4540 175 176 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.n17a 175 170 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.n0 4540 4540 161 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b2.n4b 4540 163 164 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b2.n16a 170 4478 201 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_b2.n16b 201 4478 170 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_b2.n15c 177 4535 201 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b2.n17b 4540 170 175 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.n18a 176 175 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.n6d 167 164 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b2.n3 162 161 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b2.n7d 4541 171 200 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b2.n5a 171 162 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b2.n7c 200 171 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b2.n18e 176 175 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.n6c 4541 164 167 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b2.n14b 201 200 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b2.n6b 167 164 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b2.n7b 4541 171 200 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b2.n15a 177 4535 201 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b2.n7a 200 171 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b2.n6a 4541 164 167 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b2.n8d 167 4535 166 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b2.n8c 166 4535 167 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b2.n8b 167 4535 166 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b2.n8a 166 4535 167 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b2.n18b 4540 175 176 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.n4a 164 163 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b2.n17c 175 170 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b2.n14c 4541 200 201 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b2.n15d 201 4535 177 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b2.n2 162 4540 163 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b2.n5b 4540 162 171 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b2.n18c 176 175 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.n17d 4540 509 475 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.n14a 4541 686 508 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_noe.n18f 4540 475 431 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.n16c 509 4478 508 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_noe.n15b 508 4535 738 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_noe.n1 4540 4540 739 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_noe.n14d 508 686 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_noe.n16d 508 4478 509 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_noe.n18d 4540 475 431 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.n17a 475 509 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.n0 4540 4540 688 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_noe.n4b 4540 687 684 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_noe.n16a 509 4478 508 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_noe.n16b 508 4478 509 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_noe.n15c 738 4535 508 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_noe.n17b 4540 509 475 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.n18a 431 475 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.n6d 685 684 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_noe.n3 739 688 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_noe.n7d 4541 740 686 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_noe.n5a 740 739 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_noe.n7c 686 740 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_noe.n18e 431 475 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.n6c 4541 684 685 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_noe.n14b 508 686 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_noe.n6b 685 684 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_noe.n7b 4541 740 686 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_noe.n15a 738 4535 508 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_noe.n7a 686 740 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_noe.n6a 4541 684 685 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_noe.n8d 685 4535 736 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_noe.n8c 736 4535 685 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_noe.n8b 685 4535 736 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_noe.n8a 736 4535 685 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_noe.n18b 4540 475 431 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.n4a 684 687 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_noe.n17c 475 509 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_noe.n14c 4541 686 508 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_noe.n15d 508 4535 738 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_noe.n2 739 4540 687 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_noe.n5b 4540 739 740 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_noe.n18c 431 475 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.n16b 4540 4478 3408 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_ng.n1 4540 3493 3576 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_ng.n17a 3407 3408 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.n18d 4540 3407 3235 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.n14d 3301 3456 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ng.n16d 4540 4478 3408 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_ng.n16a 3408 4478 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_ng.n15b 3301 4535 3573 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ng.n14a 4541 3456 3301 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ng.n16c 3408 4478 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_ng.n18f 4540 3407 3235 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.n18c 3235 3407 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.n17d 4540 3408 3407 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.n5b 4540 3576 3575 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_ng.n14c 4541 3456 3301 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ng.n2 3576 4478 3574 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_ng.n15d 3301 4535 3573 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ng.n18b 4540 3407 3235 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.n17c 3407 3408 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.n8a 3663 4535 3455 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ng.n8b 3455 4535 3663 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ng.n8c 3663 4535 3455 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ng.n8d 3455 4535 3663 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ng.n6a 4541 3457 3455 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ng.n14b 3301 3456 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ng.n7a 3456 3575 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ng.n15a 3573 4535 3301 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ng.n4a 3457 3574 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_ng.n5a 3575 3576 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_ng.n7b 4541 3575 3456 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ng.n3 3576 3577 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_ng.n6b 3455 3457 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ng.n6c 4541 3457 3455 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ng.n18a 3235 3407 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.n7c 3456 3575 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ng.n18e 3235 3407 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.n7d 4541 3575 3456 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ng.n17b 4540 3408 3407 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_ng.n6d 3455 3457 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_ng.n15c 3573 4535 3301 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_ng.n4b 4540 3574 3457 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_ng.n0 4540 4478 3577 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i0.n17d 4540 120 121 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.n14a 4541 45 119 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i0.n18f 4540 121 131 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.n16c 120 4478 119 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i0.n15b 119 4535 44 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i0.n1 4540 4540 118 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i0.n14d 119 45 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i0.n16d 119 4478 120 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i0.n18d 4540 121 131 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.n17a 121 120 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.n0 4540 4540 115 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i0.n4b 4540 116 117 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i0.n16a 120 4478 119 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i0.n16b 119 4478 120 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i0.n15c 44 4535 119 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i0.n17b 4540 120 121 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.n18a 131 121 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.n6d 43 117 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i0.n3 118 115 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i0.n7d 4541 114 45 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i0.n5a 114 118 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i0.n7c 45 114 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i0.n18e 131 121 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.n6c 4541 117 43 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i0.n14b 119 45 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i0.n6b 43 117 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i0.n7b 4541 114 45 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i0.n15a 44 4535 119 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i0.n7a 45 114 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i0.n6a 4541 117 43 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i0.n8d 43 4535 41 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i0.n8c 41 4535 43 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i0.n8b 43 4535 41 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i0.n8a 41 4535 43 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i0.n18b 4540 121 131 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.n4a 117 116 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i0.n17c 121 120 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i0.n14c 4541 45 119 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i0.n15d 119 4535 44 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i0.n2 118 4540 116 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i0.n5b 4540 118 114 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i0.n18c 131 121 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.n17d 4540 3025 3132 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.n14a 4541 3134 3135 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a1.n18f 4540 3132 3133 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.n16c 3025 4478 3135 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_a1.n15b 3135 4535 3136 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a1.n1 4540 4540 2751 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a1.n14d 3135 3134 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a1.n16d 3135 4478 3025 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_a1.n18d 4540 3132 3133 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.n17a 3132 3025 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.n0 4540 4540 2752 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a1.n4b 4540 2858 2976 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a1.n16a 3025 4478 3135 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_a1.n16b 3135 4478 3025 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_a1.n15c 3136 4535 3135 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a1.n17b 4540 3025 3132 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.n18a 3133 3132 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.n6d 2977 2976 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a1.n3 2751 2752 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a1.n7d 4541 2975 3134 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a1.n5a 2975 2751 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a1.n7c 3134 2975 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a1.n18e 3133 3132 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.n6c 4541 2976 2977 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a1.n14b 3135 3134 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a1.n6b 2977 2976 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a1.n7b 4541 2975 3134 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a1.n15a 3136 4535 3135 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a1.n7a 3134 2975 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a1.n6a 4541 2976 2977 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a1.n8d 2977 4535 2978 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a1.n8c 2978 4535 2977 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a1.n8b 2977 4535 2978 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a1.n8a 2978 4535 2977 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a1.n18b 4540 3132 3133 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.n4a 2976 2858 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a1.n17c 3132 3025 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a1.n14c 4541 3134 3135 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a1.n15d 3135 4535 3136 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a1.n2 2751 4540 2858 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a1.n5b 4540 2751 2975 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a1.n18c 3133 3132 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.n17d 4540 734 819 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.n14a 4541 821 822 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b1.n18f 4540 819 820 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.n16c 734 4478 822 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_b1.n15b 822 4535 735 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b1.n1 4540 4540 474 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b1.n14d 822 821 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b1.n16d 822 4478 734 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_b1.n18d 4540 819 820 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.n17a 819 734 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.n0 4540 4540 473 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b1.n4b 4540 506 680 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b1.n16a 734 4478 822 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_b1.n16b 822 4478 734 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_b1.n15c 735 4535 822 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b1.n17b 4540 734 819 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.n18a 820 819 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.n6d 683 680 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b1.n3 474 473 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b1.n7d 4541 681 821 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b1.n5a 681 474 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b1.n7c 821 681 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b1.n18e 820 819 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.n6c 4541 680 683 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b1.n14b 822 821 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b1.n6b 683 680 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b1.n7b 4541 681 821 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b1.n15a 735 4535 822 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b1.n7a 821 681 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b1.n6a 4541 680 683 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b1.n8d 683 4535 682 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b1.n8c 682 4535 683 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b1.n8b 683 4535 682 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b1.n8a 682 4535 683 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_b1.n18b 4540 819 820 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.n4a 680 506 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b1.n17c 819 734 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_b1.n14c 4541 821 822 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b1.n15d 822 4535 735 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_b1.n2 474 4540 506 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b1.n5b 4540 474 681 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_b1.n18c 820 819 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddick0.29onymous_ 2422 2421 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddick0.86onymous_ 2422 2121 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddick0.23onymous_ 4540 2421 2422 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddick0.81onymous_ 4540 2121 2422 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddick0.18onymous_ 2421 4476 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddick0.75onymous_ 2422 2121 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddick0.44onymous_ 2422 2421 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddick0.96onymous_ 4540 2121 2422 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddick0.70onymous_ 4540 4476 2121 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vddick0.34onymous_ 4540 2421 2422 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.n17d 4540 76 77 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.n14a 4541 20 75 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i5.n18f 4540 77 125 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.n16c 76 4478 75 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i5.n15b 75 4535 19 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i5.n1 4540 4540 71 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i5.n14d 75 20 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i5.n16d 75 4478 76 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i5.n18d 4540 77 125 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.n17a 77 76 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.n0 4540 4540 72 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i5.n4b 4540 73 74 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i5.n16a 76 4478 75 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i5.n16b 75 4478 76 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i5.n15c 19 4535 75 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i5.n17b 4540 76 77 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.n18a 125 77 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.n6d 18 74 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i5.n3 71 72 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i5.n7d 4541 70 20 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i5.n5a 70 71 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i5.n7c 20 70 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i5.n18e 125 77 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.n6c 4541 74 18 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i5.n14b 75 20 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i5.n6b 18 74 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i5.n7b 4541 70 20 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i5.n15a 19 4535 75 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i5.n7a 20 70 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i5.n6a 4541 74 18 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i5.n8d 18 4535 16 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i5.n8c 16 4535 18 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i5.n8b 18 4535 16 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i5.n8a 16 4535 18 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i5.n18b 4540 77 125 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.n4a 74 73 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i5.n17c 77 76 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i5.n14c 4541 20 75 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i5.n15d 75 4535 19 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i5.n2 71 4540 73 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i5.n5b 4540 71 70 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i5.n18c 125 77 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.n18c 4427 4426 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.n14a 4541 4503 4504 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y2.n15b 4504 4535 4537 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y2.n16c 4425 4478 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_y2.n1 4540 4423 4420 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y2.n14d 4504 4503 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y2.n18d 4540 4426 4427 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.n16d 4540 4478 4425 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_y2.n17a 4426 4425 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.n16a 4425 4478 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_y2.n4b 4540 4424 4481 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y2.n0 4540 4422 4421 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y2.n16b 4540 4478 4425 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_y2.n6d 4501 4481 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y2.n15c 4537 4535 4504 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y2.n7d 4541 4482 4503 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y2.n17b 4540 4425 4426 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.n7c 4503 4482 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y2.n4a 4481 4424 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y2.n6c 4541 4481 4501 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y2.n6b 4501 4481 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y2.n18e 4427 4426 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.n18a 4427 4426 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.n3 4420 4421 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y2.n7b 4541 4482 4503 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y2.n7a 4503 4482 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y2.n5a 4482 4420 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y2.n6a 4541 4481 4501 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y2.n15a 4537 4535 4504 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y2.n8d 4501 4535 4502 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y2.n14b 4504 4503 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y2.n8c 4502 4535 4501 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y2.n8b 4501 4535 4502 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y2.n8a 4502 4535 4501 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_y2.n17c 4426 4425 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.n2 4420 4422 4424 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y2.n18b 4540 4426 4427 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.n15d 4504 4535 4537 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y2.n18f 4540 4426 4427 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_y2.n14c 4541 4503 4504 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_y2.n5b 4540 4420 4482 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_y2.n17d 4540 4425 4426 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.n17d 4540 2466 2573 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.n14a 4541 2574 2575 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a2.n18f 4540 2573 2929 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.n16c 2466 4478 2575 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_a2.n15b 2575 4535 2467 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a2.n1 4540 4540 2243 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a2.n14d 2575 2574 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a2.n16d 2575 4478 2466 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_a2.n18d 4540 2573 2929 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.n17a 2573 2466 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.n0 4540 4540 2242 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a2.n4b 4540 2282 2417 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a2.n16a 2466 4478 2575 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_a2.n16b 2575 4478 2466 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_a2.n15c 2467 4535 2575 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a2.n17b 4540 2466 2573 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.n18a 2929 2573 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.n6d 2420 2417 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a2.n3 2243 2242 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a2.n7d 4541 2418 2574 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a2.n5a 2418 2243 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a2.n7c 2574 2418 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a2.n18e 2929 2573 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.n6c 4541 2417 2420 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a2.n14b 2575 2574 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a2.n6b 2420 2417 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a2.n7b 4541 2418 2574 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a2.n15a 2467 4535 2575 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a2.n7a 2574 2418 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a2.n6a 4541 2417 2420 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a2.n8d 2420 4535 2419 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a2.n8c 2419 4535 2420 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a2.n8b 2420 4535 2419 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a2.n8a 2419 4535 2420 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_a2.n18b 4540 2573 2929 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.n4a 2417 2282 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a2.n17c 2573 2466 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_a2.n14c 4541 2574 2575 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a2.n15d 2575 4535 2467 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_a2.n2 2243 4540 2282 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a2.n5b 4540 2243 2418 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_a2.n18c 2929 2573 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.n17d 4540 4450 4451 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.n14a 4541 4518 4519 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d3.n18f 4540 4451 4452 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.n16c 4450 4478 4519 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_d3.n15b 4519 4535 4542 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d3.n1 4540 4540 4447 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d3.n14d 4519 4518 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d3.n16d 4519 4478 4450 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_d3.n18d 4540 4451 4452 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.n17a 4451 4450 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.n0 4540 4540 4448 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d3.n4b 4540 4449 4488 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d3.n16a 4450 4478 4519 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_d3.n16b 4519 4478 4450 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_d3.n15c 4542 4535 4519 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d3.n17b 4540 4450 4451 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.n18a 4452 4451 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.n6d 4517 4488 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d3.n3 4447 4448 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d3.n7d 4541 4487 4518 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d3.n5a 4487 4447 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d3.n7c 4518 4487 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d3.n18e 4452 4451 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.n6c 4541 4488 4517 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d3.n14b 4519 4518 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d3.n6b 4517 4488 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d3.n7b 4541 4487 4518 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d3.n15a 4542 4535 4519 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d3.n7a 4518 4487 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d3.n6a 4541 4488 4517 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d3.n8d 4517 4535 4516 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d3.n8c 4516 4535 4517 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d3.n8b 4517 4535 4516 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d3.n8a 4516 4535 4517 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_d3.n18b 4540 4451 4452 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.n4a 4488 4449 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d3.n17c 4451 4450 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_d3.n14c 4541 4518 4519 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d3.n15d 4519 4535 4542 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_d3.n2 4447 4540 4449 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d3.n5b 4540 4447 4487 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_d3.n18c 4452 4451 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.n17d 4540 112 113 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.n14a 4541 40 111 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i1.n18f 4540 113 3559 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.n16c 112 4478 111 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i1.n15b 111 4535 39 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i1.n1 4540 4540 107 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i1.n14d 111 40 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i1.n16d 111 4478 112 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i1.n18d 4540 113 3559 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.n17a 113 112 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.n0 4540 4540 108 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i1.n4b 4540 109 110 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i1.n16a 112 4478 111 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i1.n16b 111 4478 112 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i1.n15c 39 4535 111 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i1.n17b 4540 112 113 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.n18a 3559 113 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.n6d 38 110 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i1.n3 107 108 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i1.n7d 4541 106 40 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i1.n5a 106 107 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i1.n7c 40 106 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i1.n18e 3559 113 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.n6c 4541 110 38 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i1.n14b 111 40 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i1.n6b 38 110 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i1.n7b 4541 106 40 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i1.n15a 39 4535 111 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i1.n7a 40 106 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i1.n6a 4541 110 38 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i1.n8d 38 4535 36 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i1.n8c 36 4535 38 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i1.n8b 38 4535 36 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i1.n8a 36 4535 38 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i1.n18b 4540 113 3559 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.n4a 110 109 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i1.n17c 113 112 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i1.n14c 4541 40 111 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i1.n15d 111 4535 39 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i1.n2 107 4540 109 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i1.n5b 4540 107 106 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i1.n18c 3559 113 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vsseck0.75onymous_ 4540 4475 4446 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vsseck0.39onymous_ 4540 4476 4477 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vsseck0.13onymous_ 4540 4477 4446 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vsseck0.34onymous_ 4446 4477 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vsseck0.65onymous_ 4446 4475 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vsseck0.91onymous_ 4475 4476 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vsseck0.28onymous_ 4540 4477 4446 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vsseck0.86onymous_ 4540 4475 4446 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vsseck0.23onymous_ 4446 4477 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_vsseck0.80onymous_ 4446 4475 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.n16b 4540 4478 4389 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_cout.n1 4540 4397 4403 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_cout.n17a 4388 4389 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.n18d 4540 4388 4382 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.n14d 4384 4395 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_cout.n16d 4540 4478 4389 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_cout.n16a 4389 4478 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_cout.n15b 4384 4535 4400 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_cout.n14a 4541 4395 4384 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_cout.n16c 4389 4478 4540 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_cout.n18f 4540 4388 4382 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.n18c 4382 4388 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.n17d 4540 4389 4388 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.n5b 4540 4403 4402 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_cout.n14c 4541 4395 4384 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_cout.n2 4403 4478 4401 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_cout.n15d 4384 4535 4400 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_cout.n18b 4540 4388 4382 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.n17c 4388 4389 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.n8a 4399 4535 4394 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cout.n8b 4394 4535 4399 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cout.n8c 4399 4535 4394 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cout.n8d 4394 4535 4399 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cout.n6a 4541 4396 4394 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cout.n14b 4384 4395 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_cout.n7a 4395 4402 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cout.n15a 4400 4535 4384 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_cout.n4a 4396 4401 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_cout.n5a 4402 4403 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_cout.n7b 4541 4402 4395 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cout.n3 4403 4404 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_cout.n6b 4394 4396 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cout.n6c 4541 4396 4394 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cout.n18a 4382 4388 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.n7c 4395 4402 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cout.n18e 4382 4388 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.n7d 4541 4402 4395 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cout.n17b 4540 4389 4388 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cout.n6d 4394 4396 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cout.n15c 4400 4535 4384 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_cout.n4b 4540 4401 4396 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_cout.n0 4540 4478 4404 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i6.n17d 4540 68 69 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.n14a 4541 15 67 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i6.n18f 4540 69 124 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.n16c 68 4478 67 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i6.n15b 67 4535 14 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i6.n1 4540 4540 64 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i6.n14d 67 15 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i6.n16d 67 4478 68 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i6.n18d 4540 69 124 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.n17a 69 68 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.n0 4540 4540 63 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i6.n4b 4540 65 66 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i6.n16a 68 4478 67 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i6.n16b 67 4478 68 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_i6.n15c 14 4535 67 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i6.n17b 4540 68 69 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.n18a 124 69 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.n6d 13 66 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i6.n3 64 63 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i6.n7d 4541 62 15 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i6.n5a 62 64 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i6.n7c 15 62 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i6.n18e 124 69 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.n6c 4541 66 13 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i6.n14b 67 15 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i6.n6b 13 66 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i6.n7b 4541 62 15 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i6.n15a 14 4535 67 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i6.n7a 15 62 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i6.n6a 4541 66 13 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i6.n8d 13 4535 11 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i6.n8c 11 4535 13 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i6.n8b 13 4535 11 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i6.n8a 11 4535 13 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_i6.n18b 4540 69 124 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.n4a 66 65 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i6.n17c 69 68 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_i6.n14c 4541 15 67 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i6.n15d 67 4535 14 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_i6.n2 64 4540 65 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i6.n5b 4540 64 62 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_i6.n18c 124 69 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.n17d 4540 4398 4406 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.n14a 4541 4410 4411 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_cin.n18f 4540 4406 4407 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.n16c 4398 4478 4411 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_cin.n15b 4411 4535 4408 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_cin.n1 4540 4540 4385 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_cin.n14d 4411 4410 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_cin.n16d 4411 4478 4398 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_cin.n18d 4540 4406 4407 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.n17a 4406 4398 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.n0 4540 4540 4383 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_cin.n4b 4540 4386 4391 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_cin.n16a 4398 4478 4411 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_cin.n16b 4411 4478 4398 4541 tn L=0.32U W=1.3U AS=0.975P AD=0.975P PS=4.1U PD=4.1U 
Mp_cin.n15c 4408 4535 4411 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_cin.n17b 4540 4398 4406 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.n18a 4407 4406 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.n6d 4393 4391 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cin.n3 4385 4383 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_cin.n7d 4541 4390 4410 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cin.n5a 4390 4385 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_cin.n7c 4410 4390 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cin.n18e 4407 4406 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.n6c 4541 4391 4393 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cin.n14b 4411 4410 4541 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_cin.n6b 4393 4391 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cin.n7b 4541 4390 4410 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cin.n15a 4408 4535 4411 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_cin.n7a 4410 4390 4541 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cin.n6a 4541 4391 4393 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cin.n8d 4393 4535 4392 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cin.n8c 4392 4535 4393 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cin.n8b 4393 4535 4392 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cin.n8a 4392 4535 4393 4541 tn L=0.32U W=2.17U AS=1.6275P AD=1.6275P PS=5.85U PD=5.85U 
Mp_cin.n18b 4540 4406 4407 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.n4a 4391 4386 4540 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_cin.n17c 4406 4398 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
Mp_cin.n14c 4541 4410 4411 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_cin.n15d 4411 4535 4408 4541 tn L=0.35U W=20.3U AS=15.631P AD=15.631P PS=42.15U PD=42.15U 
Mp_cin.n2 4385 4540 4386 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_cin.n5b 4540 4385 4390 4541 tn L=0.32U W=1.32U AS=0.99P AD=0.99P PS=4.15U PD=4.15U 
Mp_cin.n18c 4407 4406 4540 4541 tn L=0.32U W=2.75U AS=2.0625P AD=2.0625P PS=7U PD=7U 
C4545 1 4541 2.1722e-14
C4544 2 4541 3.43699e-14
C4543 3 4541 1.75135e-14
C4542 4 4541 1.87984e-13
C4541 5 4541 1.91459e-14
C4540 6 4541 2.1722e-14
C4539 7 4541 3.43699e-14
C4538 8 4541 1.75135e-14
C4537 9 4541 1.87984e-13
C4536 10 4541 1.91459e-14
C4535 11 4541 2.1722e-14
C4534 12 4541 3.43699e-14
C4533 13 4541 1.75135e-14
C4532 14 4541 1.87984e-13
C4531 15 4541 1.91459e-14
C4530 16 4541 2.1722e-14
C4529 17 4541 3.43699e-14
C4528 18 4541 1.75135e-14
C4527 19 4541 1.87984e-13
C4526 20 4541 1.91459e-14
C4525 21 4541 2.1722e-14
C4524 22 4541 3.43699e-14
C4523 23 4541 1.75135e-14
C4522 24 4541 1.87984e-13
C4521 25 4541 1.91459e-14
C4520 26 4541 2.1722e-14
C4519 27 4541 3.43699e-14
C4518 28 4541 1.75135e-14
C4517 29 4541 1.87984e-13
C4516 30 4541 1.91459e-14
C4515 31 4541 2.1722e-14
C4514 32 4541 3.43699e-14
C4513 33 4541 1.75135e-14
C4512 34 4541 1.87984e-13
C4511 35 4541 1.91459e-14
C4510 36 4541 2.1722e-14
C4509 37 4541 3.43699e-14
C4508 38 4541 1.75135e-14
C4507 39 4541 1.87984e-13
C4506 40 4541 1.91459e-14
C4505 41 4541 2.1722e-14
C4504 42 4541 3.43699e-14
C4503 43 4541 1.75135e-14
C4502 44 4541 1.87984e-13
C4501 45 4541 1.91459e-14
C4500 46 4541 2.00607e-14
C4499 47 4541 7.19482e-15
C4498 48 4541 4.46878e-15
C4497 49 4541 7.37786e-15
C4496 50 4541 1.84601e-14
C4495 51 4541 5.71705e-14
C4494 52 4541 9.78565e-15
C4493 53 4541 1.57304e-14
C4492 54 4541 2.00607e-14
C4491 55 4541 4.46878e-15
C4490 56 4541 7.37786e-15
C4489 57 4541 7.19482e-15
C4488 58 4541 1.84601e-14
C4487 59 4541 5.71705e-14
C4486 60 4541 9.78565e-15
C4485 61 4541 1.57304e-14
C4484 62 4541 2.00607e-14
C4483 63 4541 4.46878e-15
C4482 64 4541 7.19482e-15
C4481 65 4541 7.37786e-15
C4480 66 4541 1.84601e-14
C4479 67 4541 5.71705e-14
C4478 68 4541 9.78565e-15
C4477 69 4541 1.57304e-14
C4476 70 4541 2.00607e-14
C4475 71 4541 7.19482e-15
C4474 72 4541 4.46878e-15
C4473 73 4541 7.37786e-15
C4472 74 4541 1.84601e-14
C4471 75 4541 5.71705e-14
C4470 76 4541 9.78565e-15
C4469 77 4541 1.57304e-14
C4468 78 4541 8.10579e-15
C4467 79 4541 8.10579e-15
C4466 80 4541 8.10579e-15
C4465 81 4541 8.10579e-15
C4464 82 4541 2.00607e-14
C4463 83 4541 7.19482e-15
C4462 84 4541 4.46878e-15
C4461 85 4541 7.37786e-15
C4460 86 4541 1.84601e-14
C4459 87 4541 5.71705e-14
C4458 88 4541 9.78565e-15
C4457 89 4541 1.57304e-14
C4456 90 4541 2.00607e-14
C4455 91 4541 4.46878e-15
C4454 92 4541 1.84601e-14
C4453 93 4541 7.37786e-15
C4452 94 4541 7.19482e-15
C4451 95 4541 5.71705e-14
C4450 96 4541 9.78565e-15
C4449 97 4541 1.57304e-14
C4448 98 4541 2.00607e-14
C4447 99 4541 4.46878e-15
C4446 100 4541 7.19482e-15
C4445 101 4541 7.37786e-15
C4444 102 4541 1.84601e-14
C4443 103 4541 5.71705e-14
C4442 104 4541 9.78565e-15
C4441 105 4541 1.57304e-14
C4440 106 4541 2.00607e-14
C4439 107 4541 7.19482e-15
C4438 108 4541 4.46878e-15
C4437 109 4541 7.37786e-15
C4436 110 4541 1.84601e-14
C4435 111 4541 5.71705e-14
C4434 112 4541 9.78565e-15
C4433 113 4541 1.57304e-14
C4432 114 4541 2.00607e-14
C4431 115 4541 4.46878e-15
C4430 116 4541 7.37786e-15
C4429 117 4541 1.84601e-14
C4428 118 4541 7.19482e-15
C4427 119 4541 5.71705e-14
C4426 120 4541 9.78565e-15
C4425 121 4541 1.57304e-14
C4424 122 4541 2.27916e-14
C4423 123 4541 1.642e-14
C4422 124 4541 2.09176e-14
C4421 125 4541 1.71696e-14
C4420 126 4541 3.45392e-14
C4419 127 4541 3.45392e-14
C4418 128 4541 2.42908e-14
C4417 129 4541 2.71061e-14
C4416 130 4541 2.15287e-14
C4415 131 4541 3.8908e-14
C4414 132 4541 1.063e-14
C4413 133 4541 7.19482e-15
C4412 134 4541 4.46878e-15
C4411 135 4541 4.77843e-14
C4410 136 4541 1.57304e-14
C4409 137 4541 7.37786e-15
C4408 138 4541 3.43699e-14
C4407 139 4541 9.78565e-15
C4406 140 4541 2.00607e-14
C4405 141 4541 1.84602e-14
C4404 142 4541 1.75135e-14
C4403 143 4541 2.1722e-14
C4402 144 4541 1.84601e-14
C4401 145 4541 1.75135e-14
C4400 146 4541 1.91459e-14
C4399 147 4541 7.37786e-15
C4398 148 4541 8.42009e-15
C4397 149 4541 9.78565e-15
C4396 150 4541 2.1722e-14
C4395 151 4541 1.77803e-13
C4394 152 4541 7.19482e-15
C4393 153 4541 4.46878e-15
C4392 154 4541 2.00607e-14
C4391 155 4541 1.57304e-14
C4390 156 4541 2.10378e-14
C4389 157 4541 1.91459e-14
C4388 158 4541 5.71705e-14
C4387 159 4541 1.87984e-13
C4386 160 4541 3.43699e-14
C4385 161 4541 4.46878e-15
C4384 162 4541 7.19482e-15
C4383 163 4541 7.37786e-15
C4382 164 4541 1.84602e-14
C4381 165 4541 3.43699e-14
C4380 166 4541 2.1722e-14
C4379 167 4541 1.75135e-14
C4378 168 4541 1.75135e-14
C4377 169 4541 1.91459e-14
C4376 170 4541 9.78565e-15
C4375 171 4541 2.00607e-14
C4374 172 4541 1.70727e-14
C4373 173 4541 5.90616e-14
C4372 174 4541 9.78565e-15
C4371 175 4541 1.57304e-14
C4370 176 4541 3.49053e-14
C4369 177 4541 1.87984e-13
C4368 178 4541 2.1722e-14
C4367 179 4541 3.43699e-14
C4366 180 4541 1.77803e-13
C4346 200 4541 1.91459e-14
C4345 201 4541 5.71705e-14
C4340 206 4541 4.48681e-15
C4339 207 4541 1.76037e-14
C4337 209 4541 4.45761e-15
C4336 210 4541 1.0065e-14
C4335 211 4541 1.1306e-14
C4334 212 4541 1.58238e-14
C4333 213 4541 7.73042e-15
C4330 216 4541 4.48681e-15
C4326 220 4541 4.45761e-15
C4324 222 4541 4.48681e-15
C4322 224 4541 5.18895e-15
C4319 227 4541 6.16744e-15
C4317 229 4541 1.67174e-14
C4315 231 4541 4.45761e-15
C4311 235 4541 4.48681e-15
C4308 238 4541 2.56359e-14
C4305 241 4541 4.45761e-15
C4301 245 4541 6.207e-15
C4299 247 4541 4.66356e-15
C4298 248 4541 6.53092e-15
C4297 249 4541 6.47294e-15
C4296 250 4541 1.19344e-14
C4295 251 4541 5.50197e-15
C4294 252 4541 1.11718e-15
C4293 253 4541 1.0971e-14
C4291 255 4541 1.8319e-14
C4289 257 4541 4.49173e-15
C4288 258 4541 1.28168e-14
C4287 259 4541 1.12063e-15
C4283 263 4541 4.48681e-15
C4282 264 4541 5.58114e-14
C4281 265 4541 3.57168e-14
C4279 267 4541 4.45761e-15
C4275 271 4541 6.53092e-15
C4274 272 4541 4.66356e-15
C4272 274 4541 5.50197e-15
C4271 275 4541 6.207e-15
C4269 277 4541 6.47294e-15
C4268 278 4541 1.19344e-14
C4267 279 4541 1.11718e-15
C4266 280 4541 1.0971e-14
C4263 283 4541 1.28168e-14
C4262 284 4541 4.49173e-15
C4261 285 4541 1.12063e-15
C4258 288 4541 1.25479e-14
C4256 290 4541 4.48681e-15
C4255 291 4541 3.62246e-14
C4252 294 4541 4.48681e-15
C4250 296 4541 2.09554e-14
C4246 300 4541 1.34777e-14
C4244 302 4541 4.45761e-15
C4243 303 4541 3.18208e-14
C4242 304 4541 4.45761e-15
C4240 306 4541 1.12063e-15
C4237 309 4541 4.66281e-15
C4236 310 4541 6.54238e-15
C4234 312 4541 6.21252e-15
C4232 314 4541 6.48499e-15
C4231 315 4541 5.5213e-15
C4229 317 4541 1.09972e-14
C4226 320 4541 1.30812e-14
C4225 321 4541 1.19753e-14
C4222 324 4541 1.12063e-15
C4221 325 4541 4.49173e-15
C4220 326 4541 1.27666e-14
C4218 328 4541 2.94323e-14
C4214 332 4541 3.64465e-14
C4213 333 4541 1.11718e-15
C4211 335 4541 1.39227e-14
C4210 336 4541 4.50098e-15
C4209 337 4541 1.12063e-15
C4208 338 4541 1.11718e-15
C4205 341 4541 6.53092e-15
C4204 342 4541 1.5834e-14
C4203 343 4541 4.66356e-15
C4198 348 4541 6.207e-15
C4197 349 4541 6.47294e-15
C4196 350 4541 1.0971e-14
C4195 351 4541 1.19344e-14
C4194 352 4541 5.50197e-15
C4193 353 4541 6.54238e-15
C4190 356 4541 4.66281e-15
C4188 358 4541 6.21252e-15
C4187 359 4541 6.48499e-15
C4186 360 4541 1.19753e-14
C4185 361 4541 5.5213e-15
C4184 362 4541 1.09972e-14
C4183 363 4541 5.56405e-15
C4181 365 4541 2.19632e-14
C4179 367 4541 1.52277e-14
C4177 369 4541 6.53092e-15
C4176 370 4541 4.66356e-15
C4174 372 4541 5.50197e-15
C4172 374 4541 6.207e-15
C4171 375 4541 1.39602e-14
C4170 376 4541 6.47294e-15
C4169 377 4541 1.0971e-14
C4168 378 4541 1.19344e-14
C4167 379 4541 1.6775e-15
C4166 380 4541 1.1838e-14
C4165 381 4541 9.72234e-15
C4164 382 4541 4.48681e-15
C4163 383 4541 7.15239e-15
C4162 384 4541 4.48681e-15
C4161 385 4541 1.99364e-14
C4160 386 4541 4.48681e-15
C4158 388 4541 6.53092e-15
C4157 389 4541 4.66356e-15
C4155 391 4541 6.207e-15
C4154 392 4541 6.47294e-15
C4153 393 4541 5.50197e-15
C4151 395 4541 1.0971e-14
C4150 396 4541 1.19344e-14
C4149 397 4541 1.25918e-14
C4148 398 4541 4.50098e-15
C4146 400 4541 1.2536e-14
C4145 401 4541 2.02127e-14
C4144 402 4541 1.79336e-14
C4143 403 4541 4.48681e-15
C4142 404 4541 1.8799e-14
C4141 405 4541 4.48681e-15
C4140 406 4541 3.5213e-14
C4139 407 4541 5.48163e-15
C4138 408 4541 4.48681e-15
C4137 409 4541 1.20738e-14
C4136 410 4541 4.50098e-15
C4134 412 4541 4.66281e-15
C4131 415 4541 6.54238e-15
C4130 416 4541 1.56352e-14
C4129 417 4541 1.09972e-14
C4128 418 4541 5.5213e-15
C4126 420 4541 6.21252e-15
C4125 421 4541 6.48499e-15
C4124 422 4541 1.19753e-14
C4123 423 4541 4.45761e-15
C4122 424 4541 6.53092e-15
C4120 426 4541 4.66356e-15
C4118 428 4541 6.207e-15
C4117 429 4541 5.50197e-15
C4115 431 4541 6.52028e-14
C4114 432 4541 6.47294e-15
C4113 433 4541 1.19344e-14
C4112 434 4541 1.0971e-14
C4111 435 4541 1.28168e-14
C4110 436 4541 4.49173e-15
C4108 438 4541 6.98083e-15
C4107 439 4541 4.48681e-15
C4106 440 4541 1.41505e-14
C4105 441 4541 1.9305e-14
C4102 444 4541 6.54238e-15
C4101 445 4541 4.66281e-15
C4099 447 4541 6.21252e-15
C4098 448 4541 6.48499e-15
C4097 449 4541 1.19753e-14
C4096 450 4541 5.5213e-15
C4095 451 4541 1.09972e-14
C4094 452 4541 1.20738e-14
C4093 453 4541 4.50098e-15
C4091 455 4541 1.42457e-14
C4090 456 4541 4.03312e-15
C4088 458 4541 1.42921e-14
C4087 459 4541 5.76665e-15
C4085 461 4541 4.49173e-15
C4083 463 4541 6.53092e-15
C4082 464 4541 1.55957e-14
C4081 465 4541 4.66356e-15
C4078 468 4541 6.207e-15
C4077 469 4541 6.47294e-15
C4076 470 4541 5.50197e-15
C4075 471 4541 1.19344e-14
C4074 472 4541 1.0971e-14
C4073 473 4541 4.46878e-15
C4072 474 4541 7.19482e-15
C4071 475 4541 1.57304e-14
C4069 477 4541 2.2158e-15
C4067 479 4541 9.90628e-15
C4063 483 4541 1.94492e-15
C4040 506 4541 7.37786e-15
C4039 507 4541 3.43699e-14
C4038 508 4541 5.71705e-14
C4037 509 4541 9.78565e-15
C4036 510 4541 1.2801e-14
C4035 511 4541 1.43074e-14
C4034 512 4541 1.12063e-15
C4033 513 4541 5.7126e-15
C4031 515 4541 7.20137e-15
C4030 516 4541 1.01722e-14
C4029 517 4541 1.12063e-15
C4026 520 4541 6.82881e-15
C4025 521 4541 1.17938e-14
C4019 527 4541 6.21252e-15
C4018 528 4541 4.66281e-15
C4017 529 4541 6.54238e-15
C4015 531 4541 6.48499e-15
C4013 533 4541 5.5213e-15
C4011 535 4541 1.09972e-14
C4010 536 4541 1.19753e-14
C4009 537 4541 2.67709e-14
C4005 541 4541 1.13637e-14
C4003 543 4541 6.14336e-15
C4002 544 4541 1.81794e-14
C4001 545 4541 4.45761e-15
C3999 547 4541 1.88773e-14
C3997 549 4541 4.45761e-15
C3996 550 4541 4.50098e-15
C3993 553 4541 1.23174e-14
C3992 554 4541 1.11718e-15
C3991 555 4541 2.1975e-14
C3986 560 4541 1.12063e-15
C3985 561 4541 6.207e-15
C3983 563 4541 4.66356e-15
C3982 564 4541 6.53092e-15
C3980 566 4541 6.47294e-15
C3979 567 4541 1.19344e-14
C3978 568 4541 5.50197e-15
C3977 569 4541 1.0971e-14
C3974 572 4541 1.26748e-14
C3973 573 4541 1.25918e-14
C3972 574 4541 4.50098e-15
C3971 575 4541 1.11718e-15
C3970 576 4541 2.352e-14
C3966 580 4541 4.74346e-15
C3965 581 4541 2.8569e-14
C3963 583 4541 4.45761e-15
C3957 589 4541 6.53092e-15
C3955 591 4541 6.207e-15
C3953 593 4541 4.66356e-15
C3952 594 4541 6.47294e-15
C3949 597 4541 5.50197e-15
C3948 598 4541 1.0971e-14
C3947 599 4541 1.19344e-14
C3946 600 4541 1.28168e-14
C3945 601 4541 4.49173e-15
C3944 602 4541 1.12063e-15
C3943 603 4541 1.25479e-14
C3941 605 4541 2.87317e-14
C3938 608 4541 1.33524e-14
C3934 612 4541 4.48681e-15
C3932 614 4541 1.88581e-14
C3930 616 4541 4.66281e-15
C3929 617 4541 6.54238e-15
C3926 620 4541 5.5213e-15
C3924 622 4541 6.21252e-15
C3922 624 4541 1.09972e-14
C3921 625 4541 6.48499e-15
C3920 626 4541 1.28562e-14
C3919 627 4541 1.19753e-14
C3916 630 4541 1.66961e-14
C3915 631 4541 1.11718e-15
C3914 632 4541 4.50098e-15
C3913 633 4541 3.4972e-14
C3911 635 4541 4.45761e-15
C3909 637 4541 6.53092e-15
C3906 640 4541 4.66356e-15
C3905 641 4541 6.207e-15
C3902 644 4541 6.47294e-15
C3900 646 4541 1.0971e-14
C3899 647 4541 1.19344e-14
C3898 648 4541 5.50197e-15
C3897 649 4541 1.54205e-14
C3895 651 4541 1.28168e-14
C3893 653 4541 4.49173e-15
C3892 654 4541 1.51928e-14
C3891 655 4541 1.12063e-15
C3890 656 4541 1.12063e-15
C3889 657 4541 4.49173e-15
C3888 658 4541 3.60688e-14
C3885 661 4541 3.61215e-14
C3884 662 4541 1.48591e-14
C3882 664 4541 1.12063e-15
C3881 665 4541 4.49173e-15
C3879 667 4541 6.53092e-15
C3877 669 4541 1.55957e-14
C3876 670 4541 4.66356e-15
C3873 673 4541 6.207e-15
C3870 676 4541 6.47294e-15
C3869 677 4541 1.0971e-14
C3868 678 4541 1.19344e-14
C3867 679 4541 5.50197e-15
C3866 680 4541 1.84602e-14
C3865 681 4541 2.00607e-14
C3864 682 4541 2.1722e-14
C3863 683 4541 1.75135e-14
C3862 684 4541 1.84601e-14
C3861 685 4541 1.75135e-14
C3860 686 4541 1.91459e-14
C3859 687 4541 7.37786e-15
C3858 688 4541 4.46878e-15
C3857 689 4541 7.43722e-15
C3854 692 4541 1.02049e-14
C3853 693 4541 2.59111e-14
C3852 694 4541 1.34453e-14
C3851 695 4541 6.47294e-15
C3850 696 4541 1.07371e-14
C3848 698 4541 4.73203e-15
C3846 700 4541 6.47294e-15
C3845 701 4541 1.44244e-14
C3843 703 4541 8.46329e-15
C3842 704 4541 6.45499e-15
C3840 706 4541 1.38021e-14
C3839 707 4541 1.44661e-14
C3838 708 4541 5.40713e-14
C3837 709 4541 1.24541e-14
C3836 710 4541 1.43252e-14
C3833 713 4541 1.08598e-14
C3832 714 4541 3.87403e-14
C3831 715 4541 4.2591e-14
C3830 716 4541 1.32677e-14
C3826 720 4541 1.63601e-14
C3825 721 4541 1.18475e-14
C3824 722 4541 6.92856e-15
C3823 723 4541 4.70211e-14
C3822 724 4541 6.43318e-15
C3821 725 4541 1.90473e-14
C3820 726 4541 6.47294e-15
C3818 728 4541 2.98565e-14
C3816 730 4541 2.12044e-14
C3815 731 4541 8.40977e-15
C3813 733 4541 6.47294e-15
C3812 734 4541 9.78565e-15
C3811 735 4541 1.87984e-13
C3810 736 4541 2.1722e-14
C3809 737 4541 3.43699e-14
C3808 738 4541 1.87984e-13
C3807 739 4541 7.19482e-15
C3806 740 4541 2.00607e-14
C3805 741 4541 4.48681e-15
C3803 743 4541 1.18034e-14
C3802 744 4541 4.45761e-15
C3801 745 4541 1.08037e-14
C3798 748 4541 1.0971e-14
C3797 749 4541 1.19344e-14
C3796 750 4541 6.207e-15
C3795 751 4541 4.66356e-15
C3793 753 4541 6.53092e-15
C3791 755 4541 1.31451e-14
C3788 758 4541 5.50197e-15
C3785 761 4541 4.48681e-15
C3784 762 4541 1.6774e-15
C3783 763 4541 1.01019e-13
C3782 764 4541 4.45761e-15
C3781 765 4541 8.33582e-14
C3780 766 4541 1.0971e-14
C3779 767 4541 1.19344e-14
C3778 768 4541 6.207e-15
C3777 769 4541 4.66356e-15
C3775 771 4541 6.53092e-15
C3772 774 4541 5.50197e-15
C3771 775 4541 1.94492e-15
C3770 776 4541 4.49173e-15
C3769 777 4541 1.28168e-14
C3765 781 4541 6.16744e-15
C3764 782 4541 5.45129e-15
C3763 783 4541 6.31126e-15
C3761 785 4541 3.63598e-14
C3759 787 4541 1.0971e-14
C3758 788 4541 1.19344e-14
C3755 791 4541 6.53092e-15
C3754 792 4541 6.207e-15
C3752 794 4541 4.66356e-15
C3750 796 4541 1.3638e-14
C3749 797 4541 2.50453e-15
C3748 798 4541 1.92802e-15
C3747 799 4541 5.50197e-15
C3746 800 4541 3.17142e-15
C3743 803 4541 2.37705e-14
C3741 805 4541 4.48681e-15
C3739 807 4541 1.0971e-14
C3738 808 4541 1.19344e-14
C3737 809 4541 6.53092e-15
C3734 812 4541 4.66356e-15
C3733 813 4541 6.207e-15
C3728 818 4541 5.50197e-15
C3727 819 4541 1.57304e-14
C3726 820 4541 4.57745e-14
C3725 821 4541 1.91459e-14
C3724 822 4541 5.71705e-14
C3723 823 4541 5.35364e-15
C3722 824 4541 6.69178e-15
C3721 825 4541 1.11197e-14
C3720 826 4541 5.18333e-15
C3719 827 4541 5.99695e-15
C3718 828 4541 6.17202e-15
C3717 829 4541 2.1446e-14
C3716 830 4541 7.21095e-15
C3711 835 4541 4.66356e-15
C3710 836 4541 6.53092e-15
C3709 837 4541 6.207e-15
C3707 839 4541 6.47294e-15
C3706 840 4541 5.50197e-15
C3704 842 4541 1.0971e-14
C3703 843 4541 1.50454e-14
C3702 844 4541 1.19344e-14
C3701 845 4541 1.2046e-14
C3700 846 4541 1.16931e-14
C3698 848 4541 4.23664e-15
C3697 849 4541 4.48681e-15
C3694 852 4541 4.45761e-15
C3693 853 4541 1.03537e-13
C3691 855 4541 1.18171e-13
C3690 856 4541 3.02327e-14
C3687 859 4541 1.04827e-14
C3685 861 4541 6.53092e-15
C3684 862 4541 4.66356e-15
C3682 864 4541 6.207e-15
C3680 866 4541 6.47294e-15
C3679 867 4541 1.51044e-14
C3678 868 4541 5.50197e-15
C3677 869 4541 1.0971e-14
C3676 870 4541 1.19344e-14
C3675 871 4541 1.14928e-14
C3673 873 4541 4.48681e-15
C3672 874 4541 1.30023e-14
C3669 877 4541 5.25892e-14
C3666 880 4541 6.92856e-15
C3664 882 4541 2.17945e-14
C3662 884 4541 2.35262e-14
C3659 887 4541 1.5471e-14
C3658 888 4541 2.09062e-14
C3656 890 4541 6.16744e-15
C3654 892 4541 1.34235e-14
C3650 896 4541 2.87872e-14
C3648 898 4541 1.15656e-14
C3647 899 4541 4.45761e-15
C3646 900 4541 1.02049e-14
C3643 903 4541 8.42776e-15
C3642 904 4541 4.19735e-14
C3639 907 4541 1.32641e-14
C3638 908 4541 2.20232e-14
C3635 911 4541 5.45129e-15
C3633 913 4541 3.76946e-14
C3632 914 4541 1.16346e-14
C3629 917 4541 3.04477e-14
C3628 918 4541 4.45761e-15
C3626 920 4541 2.61497e-14
C3625 921 4541 1.55838e-14
C3622 924 4541 6.4951e-15
C3620 926 4541 3.89687e-14
C3617 929 4541 1.31898e-14
C3616 930 4541 2.84624e-14
C3614 932 4541 5.99972e-15
C3613 933 4541 1.17168e-14
C3612 934 4541 1.31684e-14
C3611 935 4541 4.49173e-15
C3610 936 4541 1.12063e-15
C3609 937 4541 1.56237e-14
C3608 938 4541 1.74535e-14
C3607 939 4541 1.11718e-15
C3606 940 4541 4.50098e-15
C3605 941 4541 6.53092e-15
C3603 943 4541 1.79116e-14
C3602 944 4541 4.66356e-15
C3601 945 4541 6.207e-15
C3598 948 4541 6.47294e-15
C3597 949 4541 5.50197e-15
C3596 950 4541 1.0971e-14
C3595 951 4541 1.19344e-14
C3594 952 4541 1.063e-14
C3559 987 4541 1.11718e-15
C3558 988 4541 9.36329e-15
C3553 993 4541 7.19482e-15
C3552 994 4541 4.46878e-15
C3551 995 4541 4.77843e-14
C3550 996 4541 1.57304e-14
C3549 997 4541 6.02337e-15
C3548 998 4541 4.48681e-15
C3546 1000 4541 1.08372e-14
C3545 1001 4541 1.39105e-14
C3544 1002 4541 7.0732e-15
C3543 1003 4541 2.0386e-15
C3542 1004 4541 1.28823e-14
C3541 1005 4541 1.94492e-15
C3539 1007 4541 1.07538e-14
C3538 1008 4541 1.2476e-14
C3537 1009 4541 3.99446e-15
C3535 1011 4541 4.66356e-15
C3534 1012 4541 6.53092e-15
C3533 1013 4541 1.88647e-14
C3532 1014 4541 1.0971e-14
C3531 1015 4541 5.50197e-15
C3530 1016 4541 6.207e-15
C3526 1020 4541 6.47294e-15
C3525 1021 4541 1.19344e-14
C3522 1024 4541 4.48681e-15
C3520 1026 4541 1.55139e-14
C3519 1027 4541 1.69808e-14
C3516 1030 4541 4.01652e-14
C3514 1032 4541 6.26171e-14
C3513 1033 4541 1.2179e-14
C3512 1034 4541 1.93056e-15
C3511 1035 4541 1.16783e-14
C3510 1036 4541 1.94492e-15
C3509 1037 4541 3.24646e-14
C3508 1038 4541 8.18526e-15
C3506 1040 4541 2.65213e-14
C3504 1042 4541 6.31126e-15
C3502 1044 4541 6.45195e-14
C3501 1045 4541 1.1002e-14
C3500 1046 4541 1.93056e-15
C3499 1047 4541 1.94492e-15
C3498 1048 4541 6.31126e-15
C3497 1049 4541 1.09683e-14
C3495 1051 4541 5.27774e-14
C3494 1052 4541 6.43318e-15
C3493 1053 4541 1.76471e-14
C3492 1054 4541 6.14336e-15
C3491 1055 4541 1.61573e-14
C3490 1056 4541 1.54016e-14
C3489 1057 4541 1.37755e-14
C3488 1058 4541 1.34417e-14
C3486 1060 4541 4.48681e-15
C3485 1061 4541 5.41229e-14
C3484 1062 4541 1.54924e-14
C3483 1063 4541 4.50702e-14
C3482 1064 4541 1.66432e-14
C3481 1065 4541 1.33002e-14
C3480 1066 4541 1.85507e-14
C3479 1067 4541 1.40178e-14
C3478 1068 4541 2.31405e-14
C3477 1069 4541 1.54905e-14
C3476 1070 4541 2.10043e-14
C3474 1072 4541 2.93619e-14
C3472 1074 4541 6.53092e-15
C3471 1075 4541 4.66356e-15
C3469 1077 4541 5.50197e-15
C3468 1078 4541 6.207e-15
C3466 1080 4541 1.0971e-14
C3465 1081 4541 6.47294e-15
C3464 1082 4541 1.3055e-14
C3463 1083 4541 1.19344e-14
C3462 1084 4541 1.51843e-14
C3461 1085 4541 4.50098e-15
C3459 1087 4541 6.31126e-15
C3458 1088 4541 1.3656e-14
C3456 1090 4541 5.56464e-14
C3455 1091 4541 3.54817e-14
C3454 1092 4541 3.2274e-14
C3453 1093 4541 1.93488e-15
C3452 1094 4541 2.50524e-15
C3451 1095 4541 3.46582e-14
C3450 1096 4541 2.59401e-14
C3449 1097 4541 3.17527e-15
C3448 1098 4541 1.31919e-14
C3445 1101 4541 2.24329e-14
C3443 1103 4541 1.49532e-14
C3442 1104 4541 7.37786e-15
C3441 1105 4541 3.43699e-14
C3440 1106 4541 9.78565e-15
C3438 1108 4541 4.48681e-15
C3436 1110 4541 6.83743e-15
C3435 1111 4541 1.76561e-14
C3431 1115 4541 4.45761e-15
C3430 1116 4541 1.2944e-14
C3429 1117 4541 9.3313e-15
C3428 1118 4541 1.40946e-14
C3424 1122 4541 6.4181e-15
C3423 1123 4541 1.54805e-14
C3420 1126 4541 2.18869e-14
C3418 1128 4541 6.54238e-15
C3417 1129 4541 4.66281e-15
C3416 1130 4541 6.21252e-15
C3413 1133 4541 1.52656e-14
C3412 1134 4541 6.48499e-15
C3411 1135 4541 5.5213e-15
C3410 1136 4541 1.09972e-14
C3409 1137 4541 1.19753e-14
C3408 1138 4541 1.68112e-14
C3407 1139 4541 4.50098e-15
C3406 1140 4541 1.11718e-15
C3403 1143 4541 1.04288e-14
C3402 1144 4541 5.99695e-15
C3401 1145 4541 9.12961e-15
C3399 1147 4541 1.42053e-14
C3398 1148 4541 4.95257e-15
C3396 1150 4541 2.28157e-14
C3395 1151 4541 1.12063e-15
C3394 1152 4541 4.34825e-14
C3392 1154 4541 6.16744e-15
C3390 1156 4541 1.35513e-14
C3388 1158 4541 1.6774e-15
C3387 1159 4541 1.32011e-14
C3386 1160 4541 5.44371e-14
C3383 1163 4541 6.16744e-15
C3382 1164 4541 8.75481e-15
C3380 1166 4541 1.29302e-14
C3379 1167 4541 1.51886e-14
C3377 1169 4541 1.37184e-14
C3376 1170 4541 3.01093e-14
C3375 1171 4541 1.6775e-15
C3374 1172 4541 6.43318e-15
C3371 1175 4541 2.22173e-14
C3370 1176 4541 1.36925e-14
C3368 1178 4541 4.48681e-15
C3367 1179 4541 1.98881e-14
C3366 1180 4541 2.97334e-14
C3362 1184 4541 2.26877e-14
C3359 1187 4541 6.16744e-15
C3358 1188 4541 1.88865e-14
C3357 1189 4541 1.33539e-14
C3354 1192 4541 1.88646e-14
C3353 1193 4541 1.17751e-14
C3350 1196 4541 1.45651e-14
C3349 1197 4541 4.48681e-15
C3348 1198 4541 6.92856e-15
C3346 1200 4541 2.77149e-14
C3345 1201 4541 4.49173e-15
C3344 1202 4541 1.12063e-15
C3342 1204 4541 6.8699e-15
C3340 1206 4541 3.70872e-14
C3339 1207 4541 1.28774e-14
C3338 1208 4541 1.92802e-15
C3337 1209 4541 2.50453e-15
C3334 1212 4541 3.17142e-15
C3332 1214 4541 2.89955e-14
C3330 1216 4541 1.17168e-14
C3329 1217 4541 1.34411e-14
C3327 1219 4541 1.24799e-14
C3325 1221 4541 1.18309e-14
C3324 1222 4541 1.70033e-14
C3321 1225 4541 1.147e-14
C3320 1226 4541 4.08589e-14
C3319 1227 4541 2.50524e-15
C3318 1228 4541 1.93488e-15
C3315 1231 4541 1.20634e-14
C3314 1232 4541 4.27013e-14
C3313 1233 4541 3.17527e-15
C3311 1235 4541 2.97496e-14
C3310 1236 4541 6.31699e-15
C3308 1238 4541 1.31937e-14
C3307 1239 4541 2.00607e-14
C3306 1240 4541 1.84602e-14
C3305 1241 4541 1.75135e-14
C3304 1242 4541 2.1722e-14
C3303 1243 4541 1.84601e-14
C3302 1244 4541 1.75135e-14
C3301 1245 4541 1.91459e-14
C3300 1246 4541 7.37786e-15
C3299 1247 4541 1.12063e-15
C3297 1249 4541 1.12063e-15
C3272 1274 4541 1.12063e-15
C3268 1278 4541 9.78565e-15
C3267 1279 4541 2.1722e-14
C3266 1280 4541 1.77803e-13
C3265 1281 4541 7.19482e-15
C3264 1282 4541 4.46878e-15
C3263 1283 4541 2.00607e-14
C3262 1284 4541 5.46412e-15
C3261 1285 4541 4.49173e-15
C3259 1287 4541 4.13397e-14
C3258 1288 4541 1.30832e-14
C3256 1290 4541 5.96714e-15
C3252 1294 4541 3.47597e-14
C3250 1296 4541 4.45761e-15
C3249 1297 4541 1.55846e-14
C3248 1298 4541 5.86632e-14
C3247 1299 4541 1.1913e-14
C3245 1301 4541 2.24387e-14
C3244 1302 4541 3.09657e-14
C3243 1303 4541 4.48681e-15
C3240 1306 4541 6.54238e-15
C3239 1307 4541 4.66281e-15
C3238 1308 4541 6.21252e-15
C3236 1310 4541 6.48499e-15
C3235 1311 4541 1.26409e-14
C3234 1312 4541 5.5213e-15
C3233 1313 4541 1.09972e-14
C3231 1315 4541 7.0825e-15
C3230 1316 4541 1.19753e-14
C3228 1318 4541 1.36027e-14
C3227 1319 4541 6.31126e-15
C3225 1321 4541 4.45761e-15
C3223 1323 4541 1.36186e-14
C3220 1326 4541 4.99173e-14
C3219 1327 4541 1.93488e-15
C3218 1328 4541 4.1202e-14
C3217 1329 4541 1.31158e-14
C3216 1330 4541 1.31842e-14
C3215 1331 4541 2.60964e-14
C3214 1332 4541 2.50524e-15
C3213 1333 4541 3.17527e-15
C3212 1334 4541 7.81046e-15
C3209 1337 4541 1.3414e-14
C3208 1338 4541 1.67317e-14
C3207 1339 4541 1.70811e-14
C3205 1341 4541 2.0737e-14
C3203 1343 4541 1.10019e-14
C3202 1344 4541 1.93109e-15
C3201 1345 4541 1.662e-14
C3200 1346 4541 1.94777e-15
C3199 1347 4541 4.55089e-14
C3198 1348 4541 4.07628e-14
C3197 1349 4541 1.57795e-14
C3196 1350 4541 1.32327e-14
C3195 1351 4541 1.52024e-14
C3194 1352 4541 1.79568e-14
C3193 1353 4541 1.34417e-14
C3191 1355 4541 4.48681e-15
C3189 1357 4541 3.38572e-14
C3188 1358 4541 4.66356e-15
C3186 1360 4541 6.207e-15
C3185 1361 4541 6.53092e-15
C3184 1362 4541 6.47294e-15
C3183 1363 4541 1.27573e-14
C3182 1364 4541 5.50197e-15
C3180 1366 4541 1.0971e-14
C3179 1367 4541 1.19344e-14
C3178 1368 4541 1.84682e-14
C3177 1369 4541 1.17015e-14
C3175 1371 4541 4.94586e-14
C3174 1372 4541 2.28122e-14
C3173 1373 4541 9.49869e-15
C3172 1374 4541 2.07787e-14
C3170 1376 4541 3.02136e-14
C3169 1377 4541 1.89055e-14
C3167 1379 4541 2.10031e-14
C3166 1380 4541 4.49173e-15
C3164 1382 4541 4.03018e-14
C3162 1384 4541 6.54238e-15
C3161 1385 4541 1.58602e-14
C3160 1386 4541 4.66281e-15
C3157 1389 4541 6.21252e-15
C3155 1391 4541 6.48499e-15
C3154 1392 4541 5.5213e-15
C3153 1393 4541 1.09972e-14
C3152 1394 4541 1.19753e-14
C3151 1395 4541 6.31126e-15
C3150 1396 4541 1.24183e-14
C3148 1398 4541 1.57304e-14
C3147 1399 4541 6.22657e-14
C3146 1400 4541 1.91459e-14
C3145 1401 4541 5.71705e-14
C3144 1402 4541 1.87984e-13
C3143 1403 4541 3.43699e-14
C3141 1405 4541 1.72861e-14
C3140 1406 4541 1.6775e-15
C3139 1407 4541 1.98128e-14
C3136 1410 4541 1.12063e-15
C3135 1411 4541 1.47663e-14
C3134 1412 4541 3.46043e-14
C3133 1413 4541 9.97922e-15
C3131 1415 4541 6.09391e-15
C3126 1420 4541 9.79415e-15
C3125 1421 4541 2.17968e-14
C3123 1423 4541 4.03452e-15
C3120 1426 4541 2.18314e-14
C3118 1428 4541 5.07308e-14
C3112 1434 4541 6.48499e-15
C3111 1435 4541 5.5213e-15
C3110 1436 4541 1.09972e-14
C3109 1437 4541 1.19753e-14
C3108 1438 4541 2.29563e-14
C3106 1440 4541 1.30812e-14
C3105 1441 4541 4.00814e-14
C3104 1442 4541 6.4951e-15
C3102 1444 4541 1.12063e-15
C3101 1445 4541 1.57039e-14
C3100 1446 4541 1.67256e-14
C3097 1449 4541 1.40212e-14
C3095 1451 4541 1.16842e-14
C3094 1452 4541 2.114e-14
C3092 1454 4541 1.17654e-14
C3089 1457 4541 4.03452e-15
C3088 1458 4541 1.15962e-14
C3086 1460 4541 1.13675e-14
C3084 1462 4541 5.49306e-15
C3081 1465 4541 4.55443e-15
C3078 1468 4541 8.2988e-15
C3076 1470 4541 4.03452e-15
C3074 1472 4541 2.64988e-14
C3072 1474 4541 1.5329e-14
C3070 1476 4541 1.12063e-15
C3068 1478 4541 1.563e-14
C3063 1483 4541 5.5213e-15
C3062 1484 4541 6.48499e-15
C3061 1485 4541 1.09972e-14
C3060 1486 4541 1.19753e-14
C3059 1487 4541 1.55938e-14
C3058 1488 4541 6.31699e-15
C3056 1490 4541 4.48681e-15
C3055 1491 4541 4.24303e-15
C3054 1492 4541 1.89939e-14
C3053 1493 4541 4.48681e-15
C3047 1499 4541 1.67359e-14
C3045 1501 4541 4.48681e-15
C3043 1503 4541 4.48681e-15
C3040 1506 4541 1.12063e-15
C3039 1507 4541 6.54238e-15
C3037 1509 4541 4.66281e-15
C3036 1510 4541 6.21252e-15
C3034 1512 4541 4.49173e-15
C3032 1514 4541 4.48681e-15
C3030 1516 4541 3.69069e-14
C3029 1517 4541 1.12063e-15
C3025 1521 4541 4.48681e-15
C3024 1522 4541 2.12511e-14
C3020 1526 4541 4.45761e-15
C3019 1527 4541 3.20313e-14
C3018 1528 4541 1.12063e-15
C3017 1529 4541 4.45761e-15
C3015 1531 4541 4.45761e-15
C3014 1532 4541 2.08057e-14
C3010 1536 4541 3.94745e-14
C3009 1537 4541 1.11718e-15
C3007 1539 4541 4.49173e-15
C3006 1540 4541 1.12063e-15
C3005 1541 4541 6.54238e-15
C3004 1542 4541 6.21252e-15
C3003 1543 4541 4.66281e-15
C2999 1547 4541 1.24499e-15
C2998 1548 4541 4.46878e-15
C2997 1549 4541 4.77843e-14
C2996 1550 4541 1.063e-14
C2995 1551 4541 7.99777e-15
C2994 1552 4541 4.97893e-14
C2993 1553 4541 5.99695e-15
C2990 1556 4541 5.93293e-15
C2989 1557 4541 7.69355e-15
C2988 1558 4541 8.91875e-15
C2987 1559 4541 4.86787e-15
C2986 1560 4541 9.8747e-15
C2985 1561 4541 6.31126e-15
C2983 1563 4541 1.81709e-14
C2982 1564 4541 1.12686e-13
C2981 1565 4541 2.50921e-14
C2980 1566 4541 4.48681e-15
C2979 1567 4541 1.94492e-15
C2978 1568 4541 4.45761e-15
C2977 1569 4541 1.97741e-14
C2976 1570 4541 4.48681e-15
C2975 1571 4541 1.15154e-14
C2974 1572 4541 6.60603e-15
C2973 1573 4541 4.45761e-15
C2971 1575 4541 4.66356e-15
C2970 1576 4541 6.53092e-15
C2969 1577 4541 5.50197e-15
C2967 1579 4541 6.207e-15
C2965 1581 4541 6.47294e-15
C2964 1582 4541 1.28168e-14
C2963 1583 4541 1.0971e-14
C2962 1584 4541 1.19344e-14
C2961 1585 4541 2.79649e-14
C2960 1586 4541 4.49173e-15
C2958 1588 4541 1.25479e-14
C2957 1589 4541 2.41397e-14
C2956 1590 4541 4.48681e-15
C2955 1591 4541 1.39556e-13
C2954 1592 4541 1.17659e-14
C2953 1593 4541 4.48681e-15
C2951 1595 4541 5.11826e-15
C2950 1596 4541 4.45761e-15
C2948 1598 4541 3.04011e-14
C2946 1600 4541 1.64644e-14
C2945 1601 4541 4.49173e-15
C2942 1604 4541 4.66356e-15
C2940 1606 4541 6.207e-15
C2939 1607 4541 6.53092e-15
C2938 1608 4541 1.55957e-14
C2937 1609 4541 6.47294e-15
C2936 1610 4541 5.50197e-15
C2934 1612 4541 1.0971e-14
C2933 1613 4541 1.19344e-14
C2931 1615 4541 4.66356e-15
C2929 1617 4541 6.53092e-15
C2928 1618 4541 5.50197e-15
C2926 1620 4541 6.207e-15
C2925 1621 4541 1.0971e-14
C2924 1622 4541 6.47294e-15
C2923 1623 4541 1.19344e-14
C2922 1624 4541 1.28168e-14
C2921 1625 4541 4.49173e-15
C2919 1627 4541 1.25479e-14
C2918 1628 4541 4.66281e-15
C2916 1630 4541 6.54238e-15
C2915 1631 4541 1.09972e-14
C2914 1632 4541 5.5213e-15
C2911 1635 4541 6.21252e-15
C2910 1636 4541 6.48499e-15
C2909 1637 4541 1.19753e-14
C2908 1638 4541 1.28562e-14
C2907 1639 4541 4.50098e-15
C2905 1641 4541 1.2536e-14
C2904 1642 4541 1.43118e-14
C2903 1643 4541 4.49173e-15
C2900 1646 4541 3.81622e-14
C2899 1647 4541 1.41902e-14
C2896 1650 4541 6.53092e-15
C2895 1651 4541 1.83747e-14
C2894 1652 4541 4.66356e-15
C2892 1654 4541 6.207e-15
C2890 1656 4541 6.47294e-15
C2889 1657 4541 5.50197e-15
C2888 1658 4541 1.19344e-14
C2887 1659 4541 1.0971e-14
C2886 1660 4541 7.19482e-15
C2885 1661 4541 7.37786e-15
C2884 1662 4541 1.57304e-14
C2883 1663 4541 9.78565e-15
C2879 1667 4541 1.6775e-15
C2873 1673 4541 1.94777e-15
C2863 1683 4541 1.92802e-15
C2862 1684 4541 2.50453e-15
C2861 1685 4541 3.17142e-15
C2857 1689 4541 1.84602e-14
C2856 1690 4541 3.43699e-14
C2855 1691 4541 2.1722e-14
C2854 1692 4541 1.75135e-14
C2853 1693 4541 1.75135e-14
C2852 1694 4541 1.91459e-14
C2851 1695 4541 1.84601e-14
C2850 1696 4541 6.09391e-15
C2849 1697 4541 1.50272e-14
C2846 1700 4541 8.93947e-15
C2845 1701 4541 6.14336e-15
C2844 1702 4541 1.35723e-14
C2842 1704 4541 3.97335e-14
C2841 1705 4541 1.41686e-14
C2840 1706 4541 1.04415e-14
C2839 1707 4541 1.12063e-15
C2838 1708 4541 1.28948e-14
C2837 1709 4541 6.8699e-15
C2836 1710 4541 2.18949e-14
C2833 1713 4541 5.48163e-15
C2832 1714 4541 4.48681e-15
C2830 1716 4541 6.53092e-15
C2828 1718 4541 1.80606e-14
C2827 1719 4541 4.66356e-15
C2824 1722 4541 5.50197e-15
C2823 1723 4541 6.207e-15
C2820 1726 4541 6.47294e-15
C2819 1727 4541 1.0971e-14
C2818 1728 4541 1.19344e-14
C2816 1730 4541 2.73761e-14
C2812 1734 4541 1.11718e-15
C2810 1736 4541 4.66281e-15
C2809 1737 4541 6.54238e-15
C2808 1738 4541 1.41874e-14
C2807 1739 4541 5.5213e-15
C2805 1741 4541 6.21252e-15
C2803 1743 4541 1.09972e-14
C2802 1744 4541 6.48499e-15
C2801 1745 4541 1.19753e-14
C2799 1747 4541 1.55249e-14
C2796 1750 4541 2.22523e-14
C2795 1751 4541 1.23174e-14
C2794 1752 4541 4.50098e-15
C2793 1753 4541 1.11718e-15
C2792 1754 4541 2.10582e-14
C2791 1755 4541 7.17056e-15
C2788 1758 4541 4.03452e-15
C2782 1764 4541 1.36732e-14
C2781 1765 4541 1.36869e-14
C2777 1769 4541 4.48681e-15
C2776 1770 4541 2.31204e-14
C2772 1774 4541 1.44661e-14
C2768 1778 4541 4.55443e-15
C2766 1780 4541 4.45761e-15
C2765 1781 4541 1.11718e-15
C2764 1782 4541 2.14152e-13
C2761 1785 4541 5.25751e-14
C2758 1788 4541 4.48681e-15
C2757 1789 4541 2.05093e-14
C2756 1790 4541 1.85263e-14
C2752 1794 4541 6.92018e-15
C2749 1797 4541 1.26112e-14
C2748 1798 4541 2.68129e-14
C2743 1803 4541 4.45761e-15
C2742 1804 4541 2.59345e-14
C2740 1806 4541 6.43318e-15
C2737 1809 4541 1.70448e-14
C2736 1810 4541 3.84913e-14
C2734 1812 4541 3.43803e-14
C2733 1813 4541 1.08817e-14
C2731 1815 4541 1.75753e-14
C2728 1818 4541 1.11718e-15
C2727 1819 4541 1.31976e-14
C2725 1821 4541 1.24799e-14
C2722 1824 4541 2.09509e-14
C2721 1825 4541 1.51705e-14
C2720 1826 4541 9.78565e-15
C2719 1827 4541 2.00607e-14
C2718 1828 4541 1.77803e-13
C2717 1829 4541 7.37786e-15
C2716 1830 4541 7.19482e-15
C2715 1831 4541 4.46878e-15
C2714 1832 4541 2.00607e-14
C2713 1833 4541 5.80893e-15
C2712 1834 4541 6.48338e-15
C2711 1835 4541 3.5684e-14
C2709 1837 4541 7.59155e-15
C2708 1838 4541 3.41166e-14
C2707 1839 4541 4.45761e-15
C2704 1842 4541 1.64494e-14
C2703 1843 4541 1.72946e-14
C2702 1844 4541 7.65097e-15
C2700 1846 4541 4.0288e-15
C2699 1847 4541 2.05042e-14
C2697 1849 4541 8.3353e-15
C2695 1851 4541 8.46329e-15
C2694 1852 4541 6.53092e-15
C2692 1854 4541 4.66356e-15
C2690 1856 4541 5.50197e-15
C2689 1857 4541 6.207e-15
C2687 1859 4541 6.47294e-15
C2686 1860 4541 1.0971e-14
C2685 1861 4541 1.19344e-14
C2684 1862 4541 2.38825e-14
C2683 1863 4541 1.23174e-14
C2681 1865 4541 1.62971e-14
C2680 1866 4541 4.50098e-15
C2678 1868 4541 4.66356e-15
C2677 1869 4541 6.53092e-15
C2676 1870 4541 1.50002e-14
C2674 1872 4541 5.50197e-15
C2672 1874 4541 6.207e-15
C2671 1875 4541 6.47294e-15
C2670 1876 4541 1.19344e-14
C2669 1877 4541 1.0971e-14
C2668 1878 4541 5.54023e-14
C2667 1879 4541 6.92018e-15
C2665 1881 4541 1.34296e-14
C2664 1882 4541 6.19446e-14
C2662 1884 4541 1.20968e-14
C2661 1885 4541 4.87406e-14
C2660 1886 4541 3.58137e-14
C2659 1887 4541 1.32072e-14
C2658 1888 4541 1.93056e-15
C2657 1889 4541 1.94492e-15
C2655 1891 4541 1.09683e-14
C2654 1892 4541 6.68606e-15
C2653 1893 4541 5.11109e-14
C2652 1894 4541 1.19487e-13
C2651 1895 4541 2.18594e-14
C2650 1896 4541 2.69343e-14
C2649 1897 4541 1.31568e-14
C2647 1899 4541 4.50098e-15
C2644 1902 4541 6.53092e-15
C2643 1903 4541 4.66356e-15
C2641 1905 4541 6.207e-15
C2640 1906 4541 1.5834e-14
C2639 1907 4541 6.47294e-15
C2638 1908 4541 5.50197e-15
C2637 1909 4541 1.19344e-14
C2636 1910 4541 1.0971e-14
C2635 1911 4541 6.18686e-14
C2633 1913 4541 7.61372e-15
C2632 1914 4541 1.14947e-14
C2631 1915 4541 3.41097e-14
C2630 1916 4541 1.92802e-15
C2629 1917 4541 2.50453e-15
C2628 1918 4541 3.17142e-15
C2627 1919 4541 5.99393e-15
C2626 1920 4541 1.31976e-14
C2624 1922 4541 7.62469e-15
C2623 1923 4541 1.24686e-14
C2621 1925 4541 1.77791e-14
C2620 1926 4541 4.50098e-15
C2618 1928 4541 3.23339e-14
C2616 1930 4541 6.53092e-15
C2615 1931 4541 1.5834e-14
C2614 1932 4541 4.66356e-15
C2611 1935 4541 6.207e-15
C2610 1936 4541 6.47294e-15
C2609 1937 4541 1.19344e-14
C2608 1938 4541 1.0971e-14
C2607 1939 4541 5.50197e-15
C2606 1940 4541 1.57304e-14
C2605 1941 4541 1.87984e-13
C2604 1942 4541 2.1722e-14
C2603 1943 4541 3.43699e-14
C2595 1951 4541 2.21519e-15
C2588 1958 4541 1.93488e-15
C2587 1959 4541 3.17527e-15
C2586 1960 4541 2.50524e-15
C2576 1970 4541 1.91459e-14
C2575 1971 4541 5.71705e-14
C2574 1972 4541 7.01821e-14
C2572 1974 4541 4.48681e-15
C2571 1975 4541 3.30401e-14
C2570 1976 4541 2.47311e-14
C2569 1977 4541 1.32134e-14
C2566 1980 4541 5.99695e-15
C2565 1981 4541 8.51952e-15
C2563 1983 4541 1.11718e-15
C2562 1984 4541 1.59933e-14
C2561 1985 4541 1.15992e-14
C2558 1988 4541 6.53092e-15
C2556 1990 4541 4.66356e-15
C2553 1993 4541 6.207e-15
C2551 1995 4541 6.47294e-15
C2550 1996 4541 1.0971e-14
C2549 1997 4541 1.19344e-14
C2548 1998 4541 5.50197e-15
C2547 1999 4541 2.13728e-14
C2546 2000 4541 1.11718e-15
C2545 2001 4541 4.33082e-15
C2544 2002 4541 1.18445e-13
C2543 2003 4541 9.67239e-15
C2542 2004 4541 2.64235e-14
C2541 2005 4541 1.33308e-14
C2540 2006 4541 1.11718e-15
C2538 2008 4541 9.95947e-15
C2535 2011 4541 5.99695e-15
C2534 2012 4541 1.26946e-14
C2532 2014 4541 1.11718e-15
C2531 2015 4541 4.50098e-15
C2530 2016 4541 4.45761e-15
C2526 2020 4541 2.03248e-14
C2525 2021 4541 4.03452e-15
C2524 2022 4541 1.96719e-14
C2523 2023 4541 4.18964e-14
C2520 2026 4541 1.29697e-14
C2519 2027 4541 5.33965e-14
C2515 2031 4541 1.12631e-14
C2514 2032 4541 1.32444e-14
C2513 2033 4541 1.2887e-14
C2512 2034 4541 3.71004e-14
C2511 2035 4541 1.44435e-14
C2506 2040 4541 6.14336e-15
C2505 2041 4541 2.88533e-14
C2504 2042 4541 3.59202e-14
C2503 2043 4541 1.36561e-14
C2502 2044 4541 1.88692e-14
C2496 2050 4541 1.25485e-14
C2492 2054 4541 6.14336e-15
C2491 2055 4541 5.70374e-14
C2488 2058 4541 1.12063e-15
C2487 2059 4541 8.41938e-15
C2482 2064 4541 1.68775e-14
C2481 2065 4541 3.61333e-14
C2480 2066 4541 1.45664e-14
C2476 2070 4541 4.03373e-14
C2472 2074 4541 1.11718e-15
C2471 2075 4541 1.87586e-14
C2470 2076 4541 1.32424e-14
C2467 2079 4541 5.45039e-15
C2465 2081 4541 3.50007e-14
C2462 2084 4541 1.35057e-14
C2459 2087 4541 1.50912e-14
C2458 2088 4541 2.64473e-14
C2455 2091 4541 5.99972e-15
C2454 2092 4541 1.79045e-14
C2452 2094 4541 1.13591e-14
C2451 2095 4541 1.11718e-15
C2450 2096 4541 2.5661e-14
C2449 2097 4541 4.49173e-15
C2448 2098 4541 1.12063e-15
C2447 2099 4541 3.34754e-14
C2445 2101 4541 4.66281e-15
C2443 2103 4541 6.21252e-15
C2442 2104 4541 6.54238e-15
C2441 2105 4541 6.48499e-15
C2440 2106 4541 1.58602e-14
C2439 2107 4541 5.5213e-15
C2438 2108 4541 1.09972e-14
C2437 2109 4541 1.12063e-15
C2435 2111 4541 1.33262e-13
C2434 2112 4541 1.19753e-14
C2432 2114 4541 4.0389e-15
C2429 2117 4541 1.69347e-14
C2428 2118 4541 2.05806e-14
C2426 2120 4541 4.45761e-15
C2425 2121 4541 8.10579e-15
C2424 2122 4541 6.71551e-15
C2423 2123 4541 4.0288e-15
C2420 2126 4541 6.21252e-15
C2418 2128 4541 6.54238e-15
C2417 2129 4541 4.66281e-15
C2416 2130 4541 1.35492e-14
C2415 2131 4541 6.48499e-15
C2414 2132 4541 5.5213e-15
C2412 2134 4541 1.09972e-14
C2411 2135 4541 1.19753e-14
C2410 2136 4541 3.59887e-14
C2409 2137 4541 4.45761e-15
C2408 2138 4541 2.22151e-14
C2407 2139 4541 1.39601e-14
C2406 2140 4541 1.20604e-14
C2405 2141 4541 4.50098e-15
C2403 2143 4541 2.08134e-14
C2400 2146 4541 6.49676e-15
C2399 2147 4541 1.26197e-14
C2398 2148 4541 5.99695e-15
C2397 2149 4541 4.66281e-15
C2395 2151 4541 6.54238e-15
C2393 2153 4541 1.26409e-14
C2392 2154 4541 1.09972e-14
C2391 2155 4541 5.5213e-15
C2389 2157 4541 6.21252e-15
C2388 2158 4541 6.48499e-15
C2387 2159 4541 1.19753e-14
C2386 2160 4541 1.40275e-14
C2385 2161 4541 3.35867e-14
C2384 2162 4541 6.16744e-15
C2381 2165 4541 1.26237e-14
C2380 2166 4541 1.43792e-14
C2379 2167 4541 1.72491e-14
C2378 2168 4541 4.26721e-14
C2377 2169 4541 1.6774e-15
C2376 2170 4541 2.13163e-14
C2375 2171 4541 7.24763e-14
C2374 2172 4541 1.77957e-14
C2373 2173 4541 1.137e-14
C2371 2175 4541 6.33389e-14
C2370 2176 4541 7.43566e-15
C2368 2178 4541 8.60515e-15
C2367 2179 4541 1.25534e-14
C2366 2180 4541 4.66281e-15
C2363 2183 4541 6.54238e-15
C2362 2184 4541 1.09972e-14
C2361 2185 4541 5.5213e-15
C2359 2187 4541 6.21252e-15
C2358 2188 4541 6.48499e-15
C2357 2189 4541 1.30812e-14
C2356 2190 4541 1.19753e-14
C2355 2191 4541 1.69067e-14
C2354 2192 4541 4.49173e-15
C2352 2194 4541 7.48075e-15
C2351 2195 4541 3.62757e-14
C2350 2196 4541 1.83568e-14
C2349 2197 4541 7.32026e-14
C2348 2198 4541 6.73115e-15
C2347 2199 4541 5.57723e-14
C2346 2200 4541 4.50098e-15
C2344 2202 4541 1.87977e-14
C2343 2203 4541 2.56813e-14
C2342 2204 4541 4.48681e-15
C2338 2208 4541 6.53092e-15
C2337 2209 4541 4.66356e-15
C2336 2210 4541 1.0971e-14
C2335 2211 4541 5.50197e-15
C2333 2213 4541 6.207e-15
C2332 2214 4541 6.47294e-15
C2331 2215 4541 1.3055e-14
C2330 2216 4541 1.19344e-14
C2329 2217 4541 6.92675e-14
C2328 2218 4541 4.50098e-15
C2326 2220 4541 6.36144e-14
C2324 2222 4541 6.63266e-14
C2323 2223 4541 1.36186e-14
C2321 2225 4541 4.49173e-15
C2320 2226 4541 5.99393e-15
C2319 2227 4541 6.23906e-14
C2317 2229 4541 6.00303e-14
C2314 2232 4541 6.53092e-15
C2313 2233 4541 1.74484e-14
C2312 2234 4541 4.66356e-15
C2309 2237 4541 6.207e-15
C2308 2238 4541 6.47294e-15
C2307 2239 4541 5.50197e-15
C2306 2240 4541 1.19344e-14
C2305 2241 4541 1.0971e-14
C2304 2242 4541 4.46878e-15
C2303 2243 4541 7.19482e-15
C2297 2249 4541 1.6775e-15
C2291 2255 4541 1.6774e-15
C2287 2259 4541 1.93109e-15
C2286 2260 4541 1.94777e-15
C2282 2264 4541 1.94492e-15
C2281 2265 4541 1.93056e-15
C2274 2272 4541 1.93488e-15
C2273 2273 4541 2.50524e-15
C2272 2274 4541 3.17527e-15
C2269 2277 4541 1.92802e-15
C2268 2278 4541 2.50453e-15
C2267 2279 4541 3.17142e-15
C2264 2282 4541 7.37786e-15
C2263 2283 4541 3.43699e-14
C2262 2284 4541 5.21737e-14
C2261 2285 4541 1.35519e-14
C2260 2286 4541 5.96714e-15
C2259 2287 4541 6.33431e-15
C2258 2288 4541 1.12063e-15
C2257 2289 4541 4.49173e-15
C2256 2290 4541 2.84693e-14
C2255 2291 4541 1.11718e-15
C2254 2292 4541 4.48681e-15
C2252 2294 4541 1.11718e-15
C2251 2295 4541 1.38126e-14
C2249 2297 4541 5.63948e-14
C2245 2301 4541 1.37398e-14
C2243 2303 4541 4.66356e-15
C2241 2305 4541 6.53092e-15
C2239 2307 4541 1.85231e-14
C2238 2308 4541 5.50197e-15
C2237 2309 4541 1.0971e-14
C2235 2311 4541 6.207e-15
C2234 2312 4541 6.47294e-15
C2233 2313 4541 1.19344e-14
C2231 2315 4541 7.19087e-14
C2229 2317 4541 1.2046e-14
C2226 2320 4541 9.95161e-15
C2225 2321 4541 1.12063e-15
C2224 2322 4541 1.48758e-14
C2223 2323 4541 3.74035e-14
C2222 2324 4541 7.06658e-15
C2221 2325 4541 1.23922e-13
C2219 2327 4541 1.16589e-14
C2218 2328 4541 1.17805e-14
C2214 2332 4541 1.20597e-14
C2212 2334 4541 8.00521e-15
C2211 2335 4541 4.7793e-14
C2209 2337 4541 5.27311e-14
C2208 2338 4541 1.36301e-14
C2205 2341 4541 1.66553e-14
C2201 2345 4541 1.35225e-14
C2200 2346 4541 1.18806e-14
C2194 2352 4541 3.24426e-14
C2193 2353 4541 4.49173e-15
C2192 2354 4541 1.12063e-15
C2191 2355 4541 1.17926e-14
C2190 2356 4541 4.86143e-14
C2189 2357 4541 8.3448e-14
C2186 2360 4541 6.09972e-14
C2183 2363 4541 4.50098e-15
C2181 2365 4541 1.11718e-15
C2180 2366 4541 1.27796e-14
C2176 2370 4541 6.54238e-15
C2174 2372 4541 1.37068e-14
C2173 2373 4541 4.66281e-15
C2172 2374 4541 5.5213e-15
C2169 2377 4541 6.21252e-15
C2168 2378 4541 6.48499e-15
C2167 2379 4541 1.09972e-14
C2166 2380 4541 1.19753e-14
C2162 2384 4541 1.55144e-14
C2158 2388 4541 1.65159e-14
C2156 2390 4541 7.8297e-14
C2155 2391 4541 7.63041e-15
C2154 2392 4541 1.27926e-14
C2153 2393 4541 1.12063e-15
C2152 2394 4541 1.48282e-14
C2151 2395 4541 7.9943e-15
C2147 2399 4541 1.58197e-14
C2145 2401 4541 1.24629e-14
C2144 2402 4541 1.17015e-14
C2142 2404 4541 1.93979e-14
C2139 2407 4541 1.11718e-15
C2136 2410 4541 7.13627e-14
C2135 2411 4541 1.08787e-14
C2132 2414 4541 4.96829e-14
C2131 2415 4541 2.93717e-14
C2130 2416 4541 1.33131e-14
C2129 2417 4541 1.84602e-14
C2128 2418 4541 2.00607e-14
C2127 2419 4541 2.1722e-14
C2126 2420 4541 1.75135e-14
C2125 2421 4541 8.10579e-15
C2124 2422 4541 3.45391e-14
C2123 2423 4541 7.95729e-14
C2122 2424 4541 2.24225e-14
C2120 2426 4541 1.19247e-14
C2119 2427 4541 6.48499e-15
C2118 2428 4541 6.47294e-15
C2117 2429 4541 6.16701e-14
C2114 2432 4541 1.25479e-14
C2111 2435 4541 5.39035e-14
C2110 2436 4541 6.46705e-15
C2109 2437 4541 2.82924e-14
C2108 2438 4541 2.20353e-14
C2107 2439 4541 1.22539e-14
C2106 2440 4541 1.38612e-14
C2103 2443 4541 3.07902e-14
C2102 2444 4541 2.30502e-14
C2101 2445 4541 2.03949e-14
C2099 2447 4541 7.80897e-14
C2098 2448 4541 7.10595e-15
C2097 2449 4541 1.04477e-14
C2096 2450 4541 2.33587e-14
C2095 2451 4541 6.48499e-15
C2093 2453 4541 1.4722e-14
C2092 2454 4541 6.48499e-15
C2091 2455 4541 5.84494e-14
C2089 2457 4541 2.63373e-14
C2087 2459 4541 1.27666e-14
C2086 2460 4541 6.43318e-15
C2084 2462 4541 1.23174e-14
C2083 2463 4541 2.22665e-14
C2081 2465 4541 6.47294e-15
C2080 2466 4541 9.78565e-15
C2079 2467 4541 1.87984e-13
C2078 2468 4541 6.31126e-15
C2075 2471 4541 1.04042e-14
C2074 2472 4541 1.75444e-14
C2073 2473 4541 2.21519e-15
C2070 2476 4541 1.10315e-14
C2069 2477 4541 1.6774e-15
C2067 2479 4541 1.44418e-14
C2065 2481 4541 4.45761e-15
C2064 2482 4541 1.6775e-15
C2063 2483 4541 9.99704e-15
C2061 2485 4541 1.09972e-14
C2060 2486 4541 1.19753e-14
C2059 2487 4541 6.21252e-15
C2058 2488 4541 7.04647e-14
C2056 2490 4541 6.54238e-15
C2055 2491 4541 4.66281e-15
C2052 2494 4541 5.5213e-15
C2049 2497 4541 3.82269e-14
C2048 2498 4541 1.0971e-14
C2047 2499 4541 1.19344e-14
C2046 2500 4541 6.207e-15
C2044 2502 4541 6.53092e-15
C2043 2503 4541 4.66356e-15
C2039 2507 4541 5.50197e-15
C2036 2510 4541 4.49173e-15
C2035 2511 4541 1.28168e-14
C2033 2513 4541 9.2757e-14
C2030 2516 4541 6.06794e-14
C2029 2517 4541 1.58012e-14
C2028 2518 4541 1.6774e-15
C2027 2519 4541 6.14336e-15
C2026 2520 4541 1.28594e-14
C2022 2524 4541 6.16744e-15
C2020 2526 4541 1.3418e-14
C2019 2527 4541 4.45761e-15
C2017 2529 4541 1.15667e-14
C2014 2532 4541 1.09972e-14
C2013 2533 4541 1.19753e-14
C2012 2534 4541 6.21252e-15
C2011 2535 4541 6.54238e-15
C2009 2537 4541 4.66281e-15
C2008 2538 4541 1.6018e-14
C2005 2541 4541 5.5213e-15
C2004 2542 4541 8.92563e-14
C2002 2544 4541 2.47246e-14
C2000 2546 4541 1.09972e-14
C1998 2548 4541 1.19753e-14
C1997 2549 4541 6.21252e-15
C1995 2551 4541 4.66281e-15
C1994 2552 4541 6.54238e-15
C1992 2554 4541 5.5213e-15
C1991 2555 4541 4.49173e-15
C1990 2556 4541 1.30812e-14
C1989 2557 4541 4.50098e-15
C1987 2559 4541 1.0971e-14
C1986 2560 4541 1.19344e-14
C1985 2561 4541 3.58661e-14
C1984 2562 4541 6.53092e-15
C1981 2565 4541 4.66356e-15
C1980 2566 4541 1.5834e-14
C1979 2567 4541 6.207e-15
C1974 2572 4541 5.50197e-15
C1973 2573 4541 1.57304e-14
C1972 2574 4541 1.91459e-14
C1971 2575 4541 5.71705e-14
C1970 2576 4541 4.27169e-15
C1969 2577 4541 1.19672e-14
C1967 2579 4541 5.71588e-15
C1966 2580 4541 1.11718e-15
C1965 2581 4541 1.34004e-14
C1964 2582 4541 1.15856e-14
C1962 2584 4541 3.58468e-14
C1961 2585 4541 7.25561e-15
C1960 2586 4541 1.11223e-14
C1959 2587 4541 1.1214e-14
C1958 2588 4541 4.48681e-15
C1957 2589 4541 2.16064e-14
C1956 2590 4541 4.48681e-15
C1954 2592 4541 1.74744e-14
C1953 2593 4541 1.14017e-14
C1952 2594 4541 1.27001e-14
C1951 2595 4541 1.11718e-15
C1950 2596 4541 1.26922e-14
C1948 2598 4541 1.31027e-14
C1946 2600 4541 2.34504e-14
C1945 2601 4541 1.19427e-14
C1944 2602 4541 1.12063e-15
C1942 2604 4541 6.53092e-15
C1941 2605 4541 4.66356e-15
C1939 2607 4541 6.207e-15
C1937 2609 4541 6.47294e-15
C1936 2610 4541 1.0971e-14
C1935 2611 4541 1.19344e-14
C1934 2612 4541 5.50197e-15
C1933 2613 4541 6.40216e-14
C1932 2614 4541 1.28168e-14
C1931 2615 4541 4.49173e-15
C1930 2616 4541 1.12063e-15
C1929 2617 4541 2.0463e-14
C1927 2619 4541 1.25479e-14
C1926 2620 4541 1.3607e-13
C1925 2621 4541 1.8534e-14
C1924 2622 4541 1.20955e-14
C1921 2625 4541 4.66356e-15
C1920 2626 4541 6.53092e-15
C1918 2628 4541 6.207e-15
C1917 2629 4541 6.47294e-15
C1916 2630 4541 1.19344e-14
C1915 2631 4541 5.50197e-15
C1913 2633 4541 1.0971e-14
C1912 2634 4541 1.28168e-14
C1911 2635 4541 4.27066e-14
C1910 2636 4541 3.84464e-14
C1909 2637 4541 1.12063e-15
C1908 2638 4541 4.49173e-15
C1907 2639 4541 1.25479e-14
C1905 2641 4541 1.56551e-14
C1903 2643 4541 3.30836e-14
C1901 2645 4541 4.66356e-15
C1900 2646 4541 6.53092e-15
C1899 2647 4541 1.72801e-14
C1898 2648 4541 1.0971e-14
C1897 2649 4541 5.50197e-15
C1895 2651 4541 6.207e-15
C1893 2653 4541 6.47294e-15
C1892 2654 4541 1.19344e-14
C1891 2655 4541 2.26572e-14
C1890 2656 4541 1.10888e-13
C1889 2657 4541 4.48681e-15
C1887 2659 4541 2.30955e-14
C1886 2660 4541 2.9379e-14
C1885 2661 4541 6.16744e-15
C1882 2664 4541 3.73247e-14
C1881 2665 4541 1.17862e-14
C1878 2668 4541 2.44714e-14
C1877 2669 4541 4.45761e-15
C1876 2670 4541 2.60433e-14
C1875 2671 4541 2.03869e-14
C1874 2672 4541 3.19679e-14
C1870 2676 4541 1.25102e-14
C1869 2677 4541 4.34137e-14
C1866 2680 4541 1.27453e-14
C1865 2681 4541 4.95387e-16
C1864 2682 4541 1.10514e-14
C1863 2683 4541 8.80256e-15
C1862 2684 4541 3.67777e-14
C1859 2687 4541 1.50383e-14
C1858 2688 4541 4.39326e-14
C1855 2691 4541 2.6886e-14
C1853 2693 4541 4.45761e-15
C1852 2694 4541 2.45271e-14
C1851 2695 4541 3.26472e-14
C1850 2696 4541 7.77385e-14
C1848 2698 4541 4.48681e-15
C1847 2699 4541 9.16164e-14
C1845 2701 4541 1.23174e-14
C1844 2702 4541 5.80566e-14
C1843 2703 4541 1.11718e-15
C1842 2704 4541 4.50098e-15
C1841 2705 4541 3.29279e-14
C1840 2706 4541 6.53092e-15
C1838 2708 4541 1.5834e-14
C1837 2709 4541 4.66356e-15
C1836 2710 4541 6.207e-15
C1833 2713 4541 6.47294e-15
C1832 2714 4541 5.50197e-15
C1831 2715 4541 1.0971e-14
C1830 2716 4541 1.19344e-14
C1829 2717 4541 1.063e-14
C1822 2724 4541 1.12063e-15
C1799 2747 4541 1.11718e-15
C1795 2751 4541 7.19482e-15
C1794 2752 4541 4.46878e-15
C1793 2753 4541 4.77843e-14
C1792 2754 4541 1.57304e-14
C1790 2756 4541 6.53092e-15
C1789 2757 4541 4.66356e-15
C1787 2759 4541 6.207e-15
C1786 2760 4541 6.47294e-15
C1785 2761 4541 1.55846e-14
C1784 2762 4541 1.19344e-14
C1783 2763 4541 5.50197e-15
C1781 2765 4541 1.0971e-14
C1780 2766 4541 5.76211e-15
C1778 2768 4541 6.21252e-15
C1775 2771 4541 6.54238e-15
C1774 2772 4541 4.66281e-15
C1773 2773 4541 6.48499e-15
C1772 2774 4541 1.64446e-14
C1771 2775 4541 5.5213e-15
C1770 2776 4541 1.09972e-14
C1769 2777 4541 1.19753e-14
C1768 2778 4541 5.94353e-14
C1767 2779 4541 5.01628e-14
C1765 2781 4541 8.92247e-14
C1764 2782 4541 8.8319e-14
C1763 2783 4541 2.12338e-14
C1761 2785 4541 1.37051e-14
C1760 2786 4541 5.76211e-15
C1756 2790 4541 6.42245e-14
C1754 2792 4541 1.25034e-14
C1752 2794 4541 5.99695e-15
C1748 2798 4541 1.6684e-14
C1747 2799 4541 6.41467e-15
C1746 2800 4541 1.98649e-14
C1745 2801 4541 4.14816e-14
C1744 2802 4541 5.50683e-14
C1743 2803 4541 1.55447e-14
C1742 2804 4541 1.18372e-14
C1741 2805 4541 4.45761e-15
C1740 2806 4541 8.90008e-14
C1739 2807 4541 2.37119e-14
C1737 2809 4541 7.77304e-14
C1735 2811 4541 2.51704e-14
C1734 2812 4541 7.91305e-14
C1732 2814 4541 7.33569e-14
C1729 2817 4541 1.74091e-14
C1728 2818 4541 4.48681e-15
C1727 2819 4541 4.01181e-15
C1726 2820 4541 4.01181e-15
C1725 2821 4541 2.63932e-14
C1723 2823 4541 2.81962e-14
C1721 2825 4541 8.30971e-14
C1720 2826 4541 4.49924e-14
C1719 2827 4541 3.50321e-14
C1718 2828 4541 6.43318e-15
C1717 2829 4541 1.22551e-14
C1716 2830 4541 3.15869e-14
C1715 2831 4541 1.33842e-14
C1714 2832 4541 1.32641e-14
C1713 2833 4541 5.45129e-15
C1712 2834 4541 2.63972e-14
C1711 2835 4541 1.4673e-14
C1710 2836 4541 3.28697e-14
C1709 2837 4541 2.12797e-14
C1708 2838 4541 4.48681e-15
C1707 2839 4541 1.17601e-14
C1706 2840 4541 1.97731e-14
C1705 2841 4541 1.03088e-13
C1704 2842 4541 1.23174e-14
C1703 2843 4541 4.50098e-15
C1702 2844 4541 6.33833e-14
C1700 2846 4541 3.79301e-14
C1698 2848 4541 6.53092e-15
C1697 2849 4541 4.66356e-15
C1696 2850 4541 1.5834e-14
C1693 2853 4541 6.207e-15
C1692 2854 4541 6.47294e-15
C1691 2855 4541 5.50197e-15
C1690 2856 4541 1.0971e-14
C1689 2857 4541 1.19344e-14
C1688 2858 4541 7.37786e-15
C1687 2859 4541 3.43699e-14
C1686 2860 4541 9.78565e-15
C1684 2862 4541 6.37148e-15
C1683 2863 4541 2.6864e-15
C1681 2865 4541 5.16123e-15
C1679 2867 4541 4.45761e-15
C1678 2868 4541 2.02879e-14
C1677 2869 4541 1.13649e-14
C1674 2872 4541 1.94777e-15
C1673 2873 4541 1.21407e-14
C1671 2875 4541 4.48681e-15
C1670 2876 4541 1.89225e-14
C1668 2878 4541 1.15973e-14
C1665 2881 4541 8.2069e-15
C1663 2883 4541 4.45761e-15
C1661 2885 4541 6.37148e-15
C1660 2886 4541 1.92686e-14
C1659 2887 4541 2.12608e-15
C1658 2888 4541 5.16123e-15
C1656 2890 4541 1.17453e-14
C1651 2895 4541 4.48681e-15
C1649 2897 4541 4.45761e-15
C1648 2898 4541 1.68925e-14
C1646 2900 4541 1.20112e-14
C1645 2901 4541 4.48681e-15
C1642 2904 4541 5.99695e-15
C1641 2905 4541 1.30746e-14
C1639 2907 4541 1.16056e-14
C1636 2910 4541 4.48681e-15
C1634 2912 4541 4.45761e-15
C1633 2913 4541 1.31782e-14
C1631 2915 4541 4.48681e-15
C1630 2916 4541 2.70259e-14
C1628 2918 4541 4.45761e-15
C1627 2919 4541 4.16326e-14
C1623 2923 4541 1.94492e-15
C1622 2924 4541 7.8303e-14
C1621 2925 4541 2.23774e-14
C1620 2926 4541 1.37385e-14
C1618 2928 4541 4.45761e-15
C1617 2929 4541 8.7293e-14
C1616 2930 4541 1.10962e-13
C1614 2932 4541 2.00507e-14
C1612 2934 4541 9.66321e-14
C1609 2937 4541 4.34321e-14
C1608 2938 4541 6.35081e-15
C1607 2939 4541 2.68308e-15
C1605 2941 4541 5.1587e-15
C1603 2943 4541 6.37148e-15
C1602 2944 4541 2.26886e-14
C1601 2945 4541 2.6864e-15
C1600 2946 4541 5.16123e-15
C1596 2950 4541 1.94777e-15
C1595 2951 4541 1.04404e-14
C1592 2954 4541 1.06943e-14
C1591 2955 4541 1.94777e-15
C1590 2956 4541 3.20508e-15
C1589 2957 4541 1.7068e-14
C1587 2959 4541 4.95741e-14
C1583 2963 4541 1.06761e-14
C1582 2964 4541 1.94492e-15
C1581 2965 4541 3.19931e-15
C1580 2966 4541 1.38443e-14
C1578 2968 4541 4.67407e-14
C1576 2970 4541 4.55443e-15
C1575 2971 4541 7.62024e-15
C1573 2973 4541 4.45761e-15
C1572 2974 4541 5.22046e-15
C1571 2975 4541 2.00607e-14
C1570 2976 4541 1.84602e-14
C1569 2977 4541 1.75135e-14
C1568 2978 4541 2.1722e-14
C1567 2979 4541 1.84601e-14
C1566 2980 4541 1.75135e-14
C1565 2981 4541 1.91459e-14
C1564 2982 4541 7.37786e-15
C1560 2986 4541 1.71034e-15
C1553 2993 4541 1.714e-15
C1540 3006 4541 1.714e-15
C1521 3025 4541 9.78565e-15
C1520 3026 4541 2.1722e-14
C1519 3027 4541 1.77803e-13
C1518 3028 4541 7.19482e-15
C1517 3029 4541 4.46878e-15
C1516 3030 4541 2.00607e-14
C1515 3031 4541 6.02337e-15
C1514 3032 4541 4.48681e-15
C1512 3034 4541 1.47058e-14
C1511 3035 4541 6.98561e-15
C1509 3037 4541 4.73275e-15
C1508 3038 4541 1.11151e-14
C1507 3039 4541 5.32888e-15
C1506 3040 4541 1.71034e-15
C1504 3042 4541 8.10769e-15
C1502 3044 4541 9.26263e-15
C1501 3045 4541 2.45831e-14
C1498 3048 4541 1.16006e-14
C1497 3049 4541 6.43318e-15
C1496 3050 4541 1.71034e-15
C1494 3052 4541 1.32193e-14
C1493 3053 4541 1.2843e-14
C1491 3055 4541 1.02411e-14
C1490 3056 4541 5.34334e-15
C1489 3057 4541 4.7281e-15
C1487 3059 4541 8.10596e-15
C1486 3060 4541 1.714e-15
C1484 3062 4541 6.15177e-15
C1483 3063 4541 1.6774e-15
C1482 3064 4541 1.68083e-14
C1481 3065 4541 1.56883e-14
C1480 3066 4541 1.37604e-14
C1479 3067 4541 2.03913e-15
C1478 3068 4541 1.94777e-15
C1477 3069 4541 7.05604e-15
C1476 3070 4541 2.74854e-14
C1475 3071 4541 4.45761e-15
C1473 3073 4541 2.35029e-14
C1472 3074 4541 1.6775e-15
C1471 3075 4541 4.0288e-15
C1469 3077 4541 1.60805e-14
C1468 3078 4541 1.79489e-14
C1465 3081 4541 5.99695e-15
C1464 3082 4541 2.6412e-14
C1463 3083 4541 1.43819e-14
C1462 3084 4541 8.55618e-15
C1461 3085 4541 1.22979e-14
C1460 3086 4541 5.34334e-15
C1459 3087 4541 4.7281e-15
C1457 3089 4541 8.10596e-15
C1455 3091 4541 4.19851e-14
C1451 3095 4541 1.714e-15
C1450 3096 4541 4.87878e-15
C1448 3098 4541 1.793e-14
C1447 3099 4541 1.714e-15
C1444 3102 4541 5.99695e-15
C1443 3103 4541 3.27623e-14
C1442 3104 4541 6.37148e-15
C1441 3105 4541 1.50773e-14
C1440 3106 4541 1.81384e-14
C1439 3107 4541 5.16123e-15
C1438 3108 4541 2.12608e-15
C1437 3109 4541 1.40105e-14
C1436 3110 4541 3.0395e-14
C1435 3111 4541 3.79743e-14
C1434 3112 4541 1.29288e-14
C1433 3113 4541 1.22237e-14
C1432 3114 4541 1.34522e-14
C1431 3115 4541 4.45761e-15
C1429 3117 4541 1.73649e-14
C1428 3118 4541 2.91974e-14
C1427 3119 4541 1.29288e-14
C1426 3120 4541 1.22237e-14
C1425 3121 4541 3.99446e-15
C1424 3122 4541 1.55159e-14
C1423 3123 4541 1.6082e-14
C1422 3124 4541 1.20455e-14
C1421 3125 4541 3.99446e-15
C1420 3126 4541 3.20508e-15
C1419 3127 4541 2.17874e-14
C1418 3128 4541 6.19425e-14
C1416 3130 4541 3.57209e-15
C1415 3131 4541 5.88761e-15
C1414 3132 4541 1.57304e-14
C1413 3133 4541 1.65402e-14
C1412 3134 4541 1.91459e-14
C1411 3135 4541 5.71705e-14
C1410 3136 4541 1.87984e-13
C1409 3137 4541 3.43699e-14
C1407 3139 4541 2.6864e-15
C1404 3142 4541 1.45826e-14
C1402 3144 4541 6.5978e-15
C1401 3145 4541 1.83665e-14
C1400 3146 4541 1.94777e-15
C1397 3149 4541 5.32888e-15
C1396 3150 4541 8.10769e-15
C1394 3152 4541 1.23234e-14
C1393 3153 4541 1.63075e-14
C1391 3155 4541 1.71034e-15
C1390 3156 4541 4.73275e-15
C1389 3157 4541 1.6775e-15
C1388 3158 4541 1.47088e-14
C1385 3161 4541 1.3352e-14
C1382 3164 4541 1.55006e-14
C1381 3165 4541 1.09057e-14
C1379 3167 4541 2.21519e-15
C1377 3169 4541 5.71588e-15
C1376 3170 4541 1.11718e-15
C1375 3171 4541 1.03373e-14
C1374 3172 4541 6.56124e-15
C1372 3174 4541 1.31187e-14
C1369 3177 4541 2.34144e-14
C1365 3181 4541 1.25981e-14
C1358 3188 4541 5.8058e-14
C1357 3189 4541 1.614e-14
C1356 3190 4541 1.22282e-14
C1353 3193 4541 1.94492e-15
C1352 3194 4541 1.28457e-14
C1351 3195 4541 5.34334e-15
C1349 3197 4541 8.10596e-15
C1346 3200 4541 1.24697e-14
C1345 3201 4541 4.7281e-15
C1344 3202 4541 1.714e-15
C1339 3207 4541 2.6864e-15
C1337 3209 4541 2.21356e-14
C1335 3211 4541 2.6864e-15
C1328 3218 4541 6.91729e-14
C1327 3219 4541 1.94492e-15
C1326 3220 4541 1.28642e-14
C1325 3221 4541 5.81664e-14
C1324 3222 4541 1.94492e-15
C1321 3225 4541 1.14888e-14
C1320 3226 4541 1.28538e-13
C1318 3228 4541 4.8851e-15
C1317 3229 4541 8.93288e-15
C1316 3230 4541 1.56878e-14
C1314 3232 4541 1.78334e-14
C1313 3233 4541 5.86786e-15
C1312 3234 4541 2.40696e-14
C1311 3235 4541 1.063e-14
C1310 3236 4541 6.37148e-15
C1309 3237 4541 5.16124e-15
C1307 3239 4541 2.04517e-14
C1304 3242 4541 1.71034e-15
C1303 3243 4541 5.85353e-15
C1300 3246 4541 1.94777e-15
C1299 3247 4541 4.24303e-15
C1298 3248 4541 1.94492e-15
C1295 3251 4541 1.12063e-15
C1293 3253 4541 2.14534e-14
C1292 3254 4541 1.21564e-14
C1291 3255 4541 4.45761e-15
C1289 3257 4541 5.96714e-15
C1288 3258 4541 1.30657e-14
C1286 3260 4541 1.16291e-14
C1285 3261 4541 4.45761e-15
C1284 3262 4541 5.82745e-15
C1280 3266 4541 1.714e-15
C1278 3268 4541 5.77421e-15
C1277 3269 4541 1.14431e-14
C1276 3270 4541 4.60228e-15
C1274 3272 4541 2.20284e-14
C1271 3275 4541 5.16124e-15
C1270 3276 4541 1.02436e-14
C1269 3277 4541 1.35971e-14
C1268 3278 4541 6.37148e-15
C1264 3282 4541 6.37148e-15
C1263 3283 4541 5.16124e-15
C1260 3286 4541 1.65573e-14
C1258 3288 4541 5.82745e-15
C1257 3289 4541 2.07848e-14
C1254 3292 4541 5.82745e-15
C1250 3296 4541 1.11718e-15
C1249 3297 4541 7.70082e-15
C1248 3298 4541 4.45761e-15
C1247 3299 4541 1.65361e-14
C1246 3300 4541 4.46878e-15
C1245 3301 4541 4.77843e-14
C1243 3303 4541 1.9929e-14
C1242 3304 4541 5.32888e-15
C1241 3305 4541 4.73275e-15
C1240 3306 4541 1.71034e-15
C1238 3308 4541 8.10769e-15
C1236 3310 4541 4.01892e-14
C1234 3312 4541 1.36706e-14
C1233 3313 4541 1.26364e-14
C1232 3314 4541 5.77421e-15
C1230 3316 4541 4.60228e-15
C1227 3319 4541 1.38638e-14
C1224 3322 4541 1.75991e-14
C1223 3323 4541 4.24303e-15
C1222 3324 4541 1.6775e-15
C1221 3325 4541 2.51563e-14
C1220 3326 4541 4.45761e-15
C1219 3327 4541 2.6631e-14
C1217 3329 4541 9.96846e-15
C1216 3330 4541 1.6774e-15
C1215 3331 4541 3.22065e-14
C1212 3334 4541 5.96714e-15
C1210 3336 4541 1.1679e-14
C1205 3341 4541 1.41371e-14
C1204 3342 4541 4.92923e-15
C1203 3343 4541 4.45761e-15
C1202 3344 4541 1.72113e-14
C1201 3345 4541 1.98487e-14
C1198 3348 4541 6.4181e-15
C1196 3350 4541 4.74346e-15
C1195 3351 4541 4.45761e-15
C1194 3352 4541 1.30937e-14
C1193 3353 4541 3.67896e-14
C1191 3355 4541 3.37353e-14
C1190 3356 4541 4.45761e-15
C1188 3358 4541 5.34334e-15
C1186 3360 4541 8.10596e-15
C1184 3362 4541 1.03752e-14
C1183 3363 4541 4.7281e-15
C1182 3364 4541 1.714e-15
C1180 3366 4541 4.45761e-15
C1179 3367 4541 4.75625e-14
C1178 3368 4541 6.35081e-15
C1177 3369 4541 5.1587e-15
C1176 3370 4541 1.36869e-14
C1175 3371 4541 2.68308e-15
C1174 3372 4541 1.59082e-14
C1173 3373 4541 6.35081e-15
C1172 3374 4541 2.68308e-15
C1171 3375 4541 5.1587e-15
C1170 3376 4541 8.9273e-15
C1169 3377 4541 5.08304e-14
C1168 3378 4541 1.29423e-14
C1167 3379 4541 1.22057e-14
C1166 3380 4541 6.16316e-14
C1165 3381 4541 1.6774e-15
C1164 3382 4541 4.24446e-15
C1163 3383 4541 6.33291e-15
C1162 3384 4541 4.45761e-15
C1160 3386 4541 1.53257e-14
C1159 3387 4541 6.16744e-15
C1158 3388 4541 4.01181e-15
C1157 3389 4541 5.9671e-14
C1156 3390 4541 5.67226e-14
C1155 3391 4541 6.51059e-14
C1153 3393 4541 3.19931e-15
C1152 3394 4541 1.15301e-14
C1150 3396 4541 1.01846e-14
C1149 3397 4541 6.61324e-14
C1148 3398 4541 5.16558e-15
C1147 3399 4541 5.3523e-15
C1145 3401 4541 5.96714e-15
C1143 3403 4541 7.20361e-15
C1142 3404 4541 1.02051e-14
C1141 3405 4541 7.19482e-15
C1140 3406 4541 7.37786e-15
C1139 3407 4541 1.57304e-14
C1138 3408 4541 9.78565e-15
C1137 3409 4541 2.6864e-15
C1132 3414 4541 2.12608e-15
C1131 3415 4541 4.95387e-16
C1130 3416 4541 1.6774e-15
C1127 3419 4541 1.12063e-15
C1123 3423 4541 2.53879e-15
C1120 3426 4541 1.12063e-15
C1115 3431 4541 3.32706e-14
C1112 3434 4541 1.94492e-15
C1110 3436 4541 2.12608e-15
C1106 3440 4541 1.94492e-15
C1105 3441 4541 2.6864e-15
C1103 3443 4541 2.68308e-15
C1101 3445 4541 1.92472e-14
C1099 3447 4541 3.15442e-14
C1096 3450 4541 2.00607e-14
C1095 3451 4541 1.84602e-14
C1094 3452 4541 3.43699e-14
C1093 3453 4541 2.1722e-14
C1092 3454 4541 1.75135e-14
C1091 3455 4541 1.75135e-14
C1090 3456 4541 1.91459e-14
C1089 3457 4541 1.84601e-14
C1088 3458 4541 6.37148e-15
C1087 3459 4541 5.16124e-15
C1086 3460 4541 1.16951e-14
C1083 3463 4541 9.11916e-15
C1080 3466 4541 4.45761e-15
C1079 3467 4541 6.14336e-15
C1078 3468 4541 1.14197e-14
C1076 3470 4541 1.26578e-14
C1073 3473 4541 1.06508e-15
C1072 3474 4541 1.12063e-15
C1071 3475 4541 6.37148e-15
C1070 3476 4541 5.16124e-15
C1069 3477 4541 8.74436e-15
C1067 3479 4541 1.18837e-14
C1065 3481 4541 1.29298e-14
C1064 3482 4541 6.00626e-15
C1060 3486 4541 1.25152e-14
C1059 3487 4541 4.49173e-15
C1058 3488 4541 1.67897e-14
C1057 3489 4541 1.20102e-14
C1054 3492 4541 2.81548e-14
C1053 3493 4541 4.5506e-14
C1052 3494 4541 1.11718e-15
C1051 3495 4541 1.53537e-14
C1050 3496 4541 1.78976e-14
C1049 3497 4541 1.11718e-15
C1048 3498 4541 5.59915e-15
C1047 3499 4541 2.63636e-14
C1045 3501 4541 3.34777e-14
C1044 3502 4541 1.59505e-14
C1043 3503 4541 6.51557e-14
C1041 3505 4541 6.44432e-15
C1040 3506 4541 1.33122e-14
C1039 3507 4541 1.49973e-14
C1038 3508 4541 1.12063e-15
C1037 3509 4541 4.78094e-14
C1036 3510 4541 4.45761e-15
C1032 3514 4541 3.46533e-14
C1031 3515 4541 5.16124e-15
C1030 3516 4541 8.36956e-15
C1026 3520 4541 6.37148e-15
C1025 3521 4541 4.3406e-14
C1021 3525 4541 6.44432e-15
C1020 3526 4541 4.00787e-14
C1017 3529 4541 4.48681e-15
C1015 3531 4541 1.0857e-14
C1014 3532 4541 5.05623e-14
C1013 3533 4541 1.11718e-15
C1012 3534 4541 6.37148e-15
C1011 3535 4541 5.16124e-15
C1009 3537 4541 6.28624e-14
C1008 3538 4541 1.91638e-14
C1004 3542 4541 6.35081e-15
C1003 3543 4541 5.1587e-15
C998 3548 4541 1.73266e-14
C996 3550 4541 4.45761e-15
C993 3553 4541 5.78173e-14
C992 3554 4541 1.97167e-14
C991 3555 4541 4.78036e-14
C989 3557 4541 1.94492e-15
C988 3558 4541 4.0389e-15
C987 3559 4541 1.11498e-13
C986 3560 4541 3.16477e-14
C985 3561 4541 1.19618e-14
C984 3562 4541 1.21282e-14
C983 3563 4541 1.31008e-14
C979 3567 4541 8.13149e-15
C978 3568 4541 5.76211e-15
C977 3569 4541 1.63643e-14
C976 3570 4541 1.93155e-14
C974 3572 4541 9.78565e-15
C973 3573 4541 1.77803e-13
C972 3574 4541 7.37786e-15
C971 3575 4541 2.00607e-14
C970 3576 4541 7.19482e-15
C969 3577 4541 4.46878e-15
C968 3578 4541 2.0865e-14
C967 3579 4541 6.37148e-15
C966 3580 4541 5.16123e-15
C965 3581 4541 2.6864e-15
C963 3583 4541 3.66738e-14
C962 3584 4541 2.12371e-14
C961 3585 4541 4.01181e-15
C960 3586 4541 7.29775e-15
C959 3587 4541 1.49654e-14
C957 3589 4541 2.43113e-15
C955 3591 4541 1.22822e-14
C954 3592 4541 2.4743e-14
C952 3594 4541 2.8614e-14
C951 3595 4541 1.09284e-14
C950 3596 4541 6.37148e-15
C949 3597 4541 5.16123e-15
C948 3598 4541 2.6864e-15
C947 3599 4541 2.52636e-14
C945 3601 4541 4.03312e-15
C944 3602 4541 1.37835e-14
C943 3603 4541 1.58371e-14
C942 3604 4541 1.18237e-14
C940 3606 4541 1.5463e-14
C938 3608 4541 1.06519e-14
C936 3610 4541 6.00626e-15
C935 3611 4541 2.26628e-14
C934 3612 4541 1.6774e-15
C933 3613 4541 1.63764e-14
C932 3614 4541 2.27298e-14
C930 3616 4541 1.16697e-14
C929 3617 4541 4.49173e-15
C927 3619 4541 7.27027e-14
C925 3621 4541 1.19273e-14
C924 3622 4541 1.47646e-14
C923 3623 4541 2.65117e-14
C922 3624 4541 1.40162e-14
C921 3625 4541 1.77563e-14
C920 3626 4541 1.03018e-14
C919 3627 4541 5.34265e-15
C918 3628 4541 6.14336e-15
C917 3629 4541 1.2935e-14
C916 3630 4541 1.5529e-14
C913 3633 4541 2.85785e-14
C912 3634 4541 1.08664e-14
C911 3635 4541 6.93401e-14
C910 3636 4541 2.17026e-14
C909 3637 4541 1.93287e-14
C908 3638 4541 6.8555e-14
C907 3639 4541 1.79843e-14
C906 3640 4541 3.99446e-15
C905 3641 4541 1.22057e-14
C904 3642 4541 2.01293e-14
C903 3643 4541 3.28719e-14
C902 3644 4541 3.99446e-15
C901 3645 4541 1.57574e-14
C900 3646 4541 3.35766e-14
C899 3647 4541 1.25453e-13
C896 3650 4541 2.38608e-14
C895 3651 4541 1.16635e-14
C894 3652 4541 7.69355e-15
C893 3653 4541 4.86787e-15
C892 3654 4541 8.91875e-15
C891 3655 4541 2.80314e-14
C890 3656 4541 3.57209e-15
C889 3657 4541 3.5765e-15
C888 3658 4541 3.79553e-14
C887 3659 4541 6.41467e-15
C886 3660 4541 1.57304e-14
C885 3661 4541 9.37292e-14
C884 3662 4541 1.87984e-13
C883 3663 4541 2.1722e-14
C882 3664 4541 3.43699e-14
C878 3668 4541 2.12608e-15
C875 3671 4541 1.94777e-15
C868 3678 4541 1.714e-15
C861 3685 4541 1.6774e-15
C860 3686 4541 1.91459e-14
C859 3687 4541 5.71705e-14
C857 3689 4541 4.48681e-15
C856 3690 4541 1.10195e-14
C855 3691 4541 1.14133e-14
C854 3692 4541 5.99695e-15
C852 3694 4541 1.93161e-14
C850 3696 4541 4.45761e-15
C848 3698 4541 4.48681e-15
C846 3700 4541 1.21009e-14
C845 3701 4541 1.49756e-14
C841 3705 4541 6.37148e-15
C838 3708 4541 1.12063e-15
C837 3709 4541 5.16124e-15
C836 3710 4541 8.12284e-14
C835 3711 4541 4.0389e-15
C834 3712 4541 7.31269e-14
C833 3713 4541 1.12063e-15
C832 3714 4541 3.13569e-14
C831 3715 4541 7.34918e-14
C830 3716 4541 1.9994e-14
C829 3717 4541 1.07206e-14
C826 3720 4541 5.85353e-15
C822 3724 4541 1.1944e-14
C820 3726 4541 1.16645e-14
C819 3727 4541 3.11218e-14
C818 3728 4541 1.12063e-15
C817 3729 4541 1.73033e-14
C814 3732 4541 1.31142e-14
C813 3733 4541 1.4924e-14
C812 3734 4541 1.11718e-15
C811 3735 4541 9.79152e-15
C810 3736 4541 6.45339e-15
C809 3737 4541 1.94777e-15
C806 3740 4541 1.30585e-14
C805 3741 4541 4.45761e-15
C804 3742 4541 1.14671e-14
C803 3743 4541 1.94492e-15
C802 3744 4541 1.3184e-14
C801 3745 4541 4.73203e-15
C799 3747 4541 4.48681e-15
C798 3748 4541 1.62988e-14
C797 3749 4541 5.34334e-15
C794 3752 4541 8.10596e-15
C792 3754 4541 4.7281e-15
C789 3757 4541 1.714e-15
C787 3759 4541 1.714e-15
C786 3760 4541 1.59664e-14
C782 3764 4541 5.45129e-15
C780 3766 4541 1.11909e-14
C775 3771 4541 1.30875e-14
C774 3772 4541 1.44441e-14
C772 3774 4541 2.74877e-14
C768 3778 4541 4.45761e-15
C766 3780 4541 1.71034e-15
C765 3781 4541 5.27209e-14
C764 3782 4541 6.45339e-15
C763 3783 4541 1.94777e-15
C762 3784 4541 1.94492e-15
C761 3785 4541 1.08382e-14
C760 3786 4541 6.34468e-14
C759 3787 4541 4.45761e-15
C756 3790 4541 3.5765e-15
C754 3792 4541 1.37723e-14
C753 3793 4541 2.78607e-14
C752 3794 4541 4.86787e-15
C751 3795 4541 8.91876e-15
C750 3796 4541 7.69355e-15
C749 3797 4541 1.77949e-14
C748 3798 4541 5.48163e-15
C747 3799 4541 1.09984e-14
C746 3800 4541 4.48681e-15
C744 3802 4541 1.02667e-14
C743 3803 4541 4.48681e-15
C742 3804 4541 1.73056e-14
C741 3805 4541 1.11718e-15
C740 3806 4541 1.24136e-14
C738 3808 4541 3.14954e-14
C737 3809 4541 4.24446e-15
C733 3813 4541 1.22226e-14
C732 3814 4541 1.33071e-14
C727 3819 4541 5.72709e-15
C726 3820 4541 5.96714e-15
C724 3822 4541 4.48681e-15
C723 3823 4541 1.56902e-14
C722 3824 4541 1.23677e-14
C721 3825 4541 1.29531e-14
C720 3826 4541 1.6774e-15
C719 3827 4541 4.24446e-15
C718 3828 4541 6.02337e-15
C717 3829 4541 3.51845e-14
C716 3830 4541 4.48681e-15
C714 3832 4541 1.01722e-14
C713 3833 4541 1.46045e-14
C711 3835 4541 1.32651e-13
C710 3836 4541 4.17877e-15
C709 3837 4541 5.71259e-15
C708 3838 4541 2.2158e-15
C707 3839 4541 3.71181e-14
C706 3840 4541 2.99129e-14
C703 3843 4541 1.19008e-14
C702 3844 4541 1.70701e-14
C700 3846 4541 8.77857e-14
C699 3847 4541 1.79586e-14
C697 3849 4541 1.6774e-15
C696 3850 4541 1.82124e-14
C695 3851 4541 1.30524e-14
C694 3852 4541 1.52452e-14
C692 3854 4541 4.49173e-15
C691 3855 4541 2.26876e-14
C690 3856 4541 4.45761e-15
C688 3858 4541 1.14682e-14
C687 3859 4541 4.48681e-15
C685 3861 4541 1.32202e-14
C684 3862 4541 4.45761e-15
C682 3864 4541 1.28824e-14
C681 3865 4541 1.39334e-14
C678 3868 4541 6.44432e-15
C677 3869 4541 4.45761e-15
C675 3871 4541 1.96971e-14
C674 3872 4541 1.2275e-14
C672 3874 4541 5.34334e-15
C671 3875 4541 4.7281e-15
C669 3877 4541 8.10596e-15
C667 3879 4541 1.714e-15
C666 3880 4541 9.46655e-15
C665 3881 4541 1.40403e-14
C664 3882 4541 4.07393e-14
C663 3883 4541 5.85353e-15
C662 3884 4541 5.28437e-15
C661 3885 4541 1.94777e-15
C660 3886 4541 1.97516e-14
C659 3887 4541 1.82276e-14
C658 3888 4541 5.32888e-15
C655 3891 4541 8.10769e-15
C653 3893 4541 4.73275e-15
C652 3894 4541 1.71034e-15
C651 3895 4541 5.78434e-15
C650 3896 4541 1.90588e-14
C647 3899 4541 6.37148e-15
C646 3900 4541 5.16123e-15
C645 3901 4541 2.12608e-15
C644 3902 4541 2.98124e-14
C643 3903 4541 3.57209e-15
C642 3904 4541 1.174e-14
C641 3905 4541 1.34518e-13
C639 3907 4541 1.53486e-14
C638 3908 4541 1.46811e-14
C636 3910 4541 3.57209e-15
C635 3911 4541 1.29028e-13
C634 3912 4541 4.48681e-15
C632 3914 4541 5.74235e-15
C631 3915 4541 1.82777e-14
C630 3916 4541 1.74038e-14
C629 3917 4541 1.24114e-14
C628 3918 4541 5.29476e-14
C626 3920 4541 6.53092e-15
C625 3921 4541 1.30209e-14
C624 3922 4541 4.66356e-15
C621 3925 4541 6.207e-15
C620 3926 4541 6.47294e-15
C619 3927 4541 5.50197e-15
C618 3928 4541 1.19344e-14
C617 3929 4541 1.0971e-14
C616 3930 4541 4.46877e-15
C615 3931 4541 4.36902e-14
C614 3932 4541 7.19482e-15
C613 3933 4541 1.57304e-14
C610 3936 4541 1.93056e-15
C609 3937 4541 2.50524e-15
C608 3938 4541 3.17527e-15
C606 3940 4541 1.6774e-15
C592 3954 4541 2.68308e-15
C590 3956 4541 1.6775e-15
C578 3968 4541 7.37786e-15
C577 3969 4541 3.43699e-14
C576 3970 4541 9.78565e-15
C575 3971 4541 5.71705e-14
C574 3972 4541 1.61327e-14
C573 3973 4541 1.51444e-14
C572 3974 4541 1.12063e-15
C569 3977 4541 1.16576e-14
C568 3978 4541 4.0389e-15
C567 3979 4541 4.48681e-15
C566 3980 4541 1.631e-14
C565 3981 4541 1.48174e-14
C564 3982 4541 1.45065e-14
C563 3983 4541 9.98149e-14
C560 3986 4541 2.93833e-14
C558 3988 4541 8.25775e-15
C556 3990 4541 1.30932e-14
C555 3991 4541 1.25813e-13
C554 3992 4541 4.45761e-15
C553 3993 4541 1.51226e-14
C552 3994 4541 3.74376e-14
C550 3996 4541 1.31633e-14
C549 3997 4541 4.24446e-15
C548 3998 4541 4.48681e-15
C547 3999 4541 8.83503e-15
C546 4000 4541 1.11718e-15
C545 4001 4541 1.25478e-14
C544 4002 4541 1.12063e-15
C543 4003 4541 1.97708e-14
C541 4005 4541 2.69603e-14
C540 4006 4541 5.96714e-15
C539 4007 4541 4.48681e-15
C538 4008 4541 1.88572e-14
C537 4009 4541 1.94492e-15
C536 4010 4541 4.05934e-14
C535 4011 4541 6.42632e-15
C533 4013 4541 4.48681e-15
C531 4015 4541 4.45761e-15
C530 4016 4541 2.598e-14
C528 4018 4541 6.45339e-15
C527 4019 4541 1.94777e-15
C526 4020 4541 1.06027e-14
C524 4022 4541 4.48681e-15
C522 4024 4541 3.84566e-14
C521 4025 4541 6.45339e-15
C520 4026 4541 1.94777e-15
C518 4028 4541 1.06027e-14
C517 4029 4541 4.48681e-15
C516 4030 4541 6.35081e-15
C514 4032 4541 4.95754e-14
C512 4034 4541 1.98329e-14
C509 4037 4541 5.1587e-15
C508 4038 4541 7.0071e-15
C507 4039 4541 3.38151e-14
C505 4041 4541 1.37249e-14
C502 4044 4541 1.2438e-14
C497 4049 4541 4.24303e-15
C495 4051 4541 1.26124e-14
C493 4053 4541 1.35541e-14
C492 4054 4541 1.48288e-14
C491 4055 4541 5.96714e-15
C490 4056 4541 1.24153e-14
C489 4057 4541 5.99695e-15
C488 4058 4541 3.74113e-14
C487 4059 4541 2.18041e-14
C485 4061 4541 5.96714e-15
C482 4064 4541 4.45761e-15
C481 4065 4541 1.87708e-14
C480 4066 4541 4.0389e-15
C479 4067 4541 1.80677e-14
C478 4068 4541 1.89003e-14
C477 4069 4541 5.99695e-15
C476 4070 4541 1.53957e-14
C475 4071 4541 9.11365e-14
C474 4072 4541 1.08761e-14
C471 4075 4541 1.84602e-14
C470 4076 4541 2.00607e-14
C469 4077 4541 2.1722e-14
C468 4078 4541 1.75135e-14
C467 4079 4541 1.84601e-14
C466 4080 4541 1.75135e-14
C465 4081 4541 1.91459e-14
C464 4082 4541 7.37786e-15
C463 4083 4541 4.46878e-15
C462 4084 4541 9.32804e-14
C458 4088 4541 6.66478e-15
C456 4090 4541 1.67992e-14
C454 4092 4541 1.192e-14
C452 4094 4541 1.59638e-14
C450 4096 4541 2.43844e-14
C448 4098 4541 2.04727e-14
C445 4101 4541 5.91127e-15
C444 4102 4541 9.39199e-14
C442 4104 4541 2.18017e-14
C441 4105 4541 1.05144e-13
C439 4107 4541 1.54082e-13
C435 4111 4541 1.95289e-14
C433 4113 4541 3.99446e-15
C431 4115 4541 6.47294e-15
C429 4117 4541 1.41072e-14
C428 4118 4541 6.48499e-15
C427 4119 4541 7.16427e-15
C425 4121 4541 7.82488e-14
C424 4122 4541 2.1578e-14
C423 4123 4541 1.2438e-14
C422 4124 4541 9.78565e-15
C421 4125 4541 1.77803e-13
C420 4126 4541 2.1722e-14
C419 4127 4541 3.43699e-14
C418 4128 4541 1.77803e-13
C417 4129 4541 7.19482e-15
C416 4130 4541 2.00607e-14
C415 4131 4541 5.96714e-15
C414 4132 4541 1.4736e-14
C412 4134 4541 5.96714e-15
C411 4135 4541 1.30026e-14
C409 4137 4541 6.36029e-14
C407 4139 4541 1.2015e-14
C405 4141 4541 6.16744e-15
C404 4142 4541 1.57621e-14
C403 4143 4541 9.11292e-15
C402 4144 4541 1.93218e-14
C400 4146 4541 3.41704e-14
C398 4148 4541 5.26427e-14
C396 4150 4541 2.6439e-14
C394 4152 4541 1.14898e-14
C392 4154 4541 4.49173e-15
C389 4157 4541 1.41021e-14
C385 4161 4541 2.35672e-14
C383 4163 4541 7.74901e-14
C382 4164 4541 1.57481e-14
C379 4167 4541 6.55542e-14
C377 4169 4541 2.79656e-14
C374 4172 4541 4.45761e-15
C373 4173 4541 5.99695e-15
C372 4174 4541 1.97282e-14
C369 4177 4541 3.53629e-14
C367 4179 4541 2.00803e-14
C366 4180 4541 4.90679e-15
C364 4182 4541 3.91998e-14
C363 4183 4541 1.6774e-15
C361 4185 4541 4.45761e-15
C360 4186 4541 3.70543e-14
C359 4187 4541 6.24015e-14
C357 4189 4541 5.16124e-15
C356 4190 4541 6.37148e-15
C355 4191 4541 1.44599e-14
C354 4192 4541 2.6864e-15
C353 4193 4541 2.6864e-15
C352 4194 4541 6.37148e-15
C351 4195 4541 5.16124e-15
C350 4196 4541 1.33456e-13
C348 4198 4541 1.25315e-13
C347 4199 4541 2.6864e-15
C344 4202 4541 1.0971e-14
C343 4203 4541 1.19344e-14
C341 4205 4541 6.53092e-15
C340 4206 4541 6.207e-15
C338 4208 4541 4.66356e-15
C336 4210 4541 1.47088e-14
C335 4211 4541 5.50197e-15
C334 4212 4541 4.45761e-15
C333 4213 4541 2.45107e-14
C332 4214 4541 4.74923e-14
C331 4215 4541 1.09972e-14
C330 4216 4541 1.19753e-14
C329 4217 4541 6.21252e-15
C327 4219 4541 4.66281e-15
C326 4220 4541 6.54238e-15
C325 4221 4541 1.59716e-14
C322 4224 4541 5.5213e-15
C321 4225 4541 1.6774e-15
C318 4228 4541 1.6774e-15
C317 4229 4541 1.57304e-14
C316 4230 4541 1.91459e-14
C315 4231 4541 5.71705e-14
C314 4232 4541 1.93787e-13
C313 4233 4541 6.77621e-14
C312 4234 4541 4.48681e-15
C311 4235 4541 7.10595e-15
C310 4236 4541 1.1935e-14
C308 4238 4541 1.78221e-14
C306 4240 4541 2.58591e-14
C305 4241 4541 2.05127e-14
C303 4243 4541 2.70897e-13
C301 4245 4541 4.45761e-15
C300 4246 4541 1.64436e-14
C299 4247 4541 1.42913e-14
C298 4248 4541 1.35592e-14
C296 4250 4541 1.02049e-14
C294 4252 4541 3.13983e-14
C293 4253 4541 2.46868e-14
C290 4256 4541 1.40352e-14
C288 4258 4541 1.91361e-14
C287 4259 4541 1.96934e-14
C286 4260 4541 1.58326e-14
C285 4261 4541 8.92018e-14
C284 4262 4541 4.21286e-14
C283 4263 4541 1.61867e-14
C282 4264 4541 1.58088e-14
C281 4265 4541 2.7759e-14
C280 4266 4541 1.49825e-14
C277 4269 4541 2.90423e-13
C276 4270 4541 1.18556e-14
C275 4271 4541 4.48681e-15
C274 4272 4541 3.78829e-14
C273 4273 4541 6.49533e-14
C271 4275 4541 1.44983e-14
C268 4278 4541 3.07305e-14
C267 4279 4541 2.25515e-14
C266 4280 4541 3.83716e-14
C265 4281 4541 4.45761e-15
C263 4283 4541 8.15627e-14
C262 4284 4541 4.11729e-14
C261 4285 4541 3.16298e-14
C260 4286 4541 5.99695e-15
C259 4287 4541 6.24179e-14
C257 4289 4541 2.30973e-14
C256 4290 4541 2.41336e-14
C254 4292 4541 2.72387e-14
C253 4293 4541 1.15534e-14
C252 4294 4541 2.96528e-14
C251 4295 4541 3.40362e-14
C250 4296 4541 1.50148e-14
C249 4297 4541 3.33104e-14
C248 4298 4541 4.42975e-14
C246 4300 4541 4.48681e-15
C245 4301 4541 5.07496e-14
C244 4302 4541 3.55969e-14
C243 4303 4541 4.11795e-14
C241 4305 4541 2.17557e-14
C239 4307 4541 6.37148e-15
C238 4308 4541 1.57889e-14
C237 4309 4541 5.16123e-15
C235 4311 4541 6.53092e-15
C234 4312 4541 4.66356e-15
C233 4313 4541 6.207e-15
C230 4316 4541 6.47294e-15
C229 4317 4541 1.19344e-14
C228 4318 4541 5.50197e-15
C227 4319 4541 1.0971e-14
C226 4320 4541 2.55811e-14
C225 4321 4541 6.58929e-15
C224 4322 4541 3.63799e-14
C222 4324 4541 1.61023e-14
C221 4325 4541 1.24202e-14
C219 4327 4541 1.59275e-14
C217 4329 4541 4.17709e-14
C215 4331 4541 5.48163e-15
C214 4332 4541 1.58392e-14
C213 4333 4541 4.48681e-15
C212 4334 4541 2.73353e-14
C210 4336 4541 4.24446e-15
C209 4337 4541 4.33883e-14
C208 4338 4541 2.54709e-14
C207 4339 4541 1.25144e-14
C206 4340 4541 4.45761e-15
C205 4341 4541 1.28736e-14
C204 4342 4541 3.73294e-14
C203 4343 4541 1.3409e-14
C202 4344 4541 1.11718e-15
C201 4345 4541 4.09669e-14
C200 4346 4541 1.24136e-14
C199 4347 4541 2.5537e-14
C197 4349 4541 4.24446e-15
C196 4350 4541 7.12469e-14
C195 4351 4541 7.22117e-14
C194 4352 4541 5.85979e-14
C193 4353 4541 4.46878e-15
C192 4354 4541 7.19482e-15
C191 4355 4541 1.57304e-14
C190 4356 4541 7.37786e-15
C189 4357 4541 3.43699e-14
C188 4358 4541 5.71705e-14
C187 4359 4541 9.78565e-15
C186 4360 4541 2.00607e-14
C185 4361 4541 1.84602e-14
C184 4362 4541 2.1722e-14
C183 4363 4541 1.75135e-14
C182 4364 4541 1.84601e-14
C181 4365 4541 1.75135e-14
C180 4366 4541 1.91459e-14
C179 4367 4541 7.37786e-15
C178 4368 4541 6.58326e-14
C177 4369 4541 9.78565e-15
C176 4370 4541 2.1722e-14
C175 4371 4541 1.77803e-13
C174 4372 4541 1.07849e-14
C173 4373 4541 7.19482e-15
C172 4374 4541 2.00607e-14
C171 4375 4541 4.46878e-15
C170 4376 4541 1.57304e-14
C169 4377 4541 8.25049e-14
C168 4378 4541 1.91459e-14
C167 4379 4541 5.71705e-14
C166 4380 4541 1.77803e-13
C165 4381 4541 3.43699e-14
C164 4382 4541 1.063e-14
C163 4383 4541 4.46878e-15
C162 4384 4541 4.77843e-14
C161 4385 4541 7.19482e-15
C160 4386 4541 7.37786e-15
C159 4387 4541 3.43699e-14
C158 4388 4541 1.57304e-14
C157 4389 4541 9.78565e-15
C156 4390 4541 2.00607e-14
C155 4391 4541 1.84602e-14
C154 4392 4541 2.1722e-14
C153 4393 4541 1.75135e-14
C152 4394 4541 1.75135e-14
C151 4395 4541 1.91459e-14
C150 4396 4541 1.84601e-14
C149 4397 4541 7.53042e-14
C148 4398 4541 9.78565e-15
C147 4399 4541 2.1722e-14
C146 4400 4541 1.77803e-13
C145 4401 4541 7.37786e-15
C144 4402 4541 2.00607e-14
C143 4403 4541 7.19482e-15
C142 4404 4541 4.46878e-15
C141 4405 4541 6.53357e-14
C140 4406 4541 1.57304e-14
C139 4407 4541 4.72737e-14
C138 4408 4541 1.87984e-13
C137 4409 4541 3.43699e-14
C136 4410 4541 1.91459e-14
C135 4411 4541 5.71705e-14
C134 4412 4541 8.54023e-15
C133 4413 4541 1.11601e-14
C132 4414 4541 7.19482e-15
C131 4415 4541 4.46878e-15
C130 4416 4541 7.37786e-15
C129 4417 4541 9.78565e-15
C128 4418 4541 1.57304e-14
C127 4419 4541 1.063e-14
C126 4420 4541 7.19482e-15
C125 4421 4541 4.46878e-15
C124 4422 4541 1.11601e-14
C123 4423 4541 8.54023e-15
C122 4424 4541 7.37786e-15
C121 4425 4541 9.78565e-15
C120 4426 4541 1.57304e-14
C119 4427 4541 1.063e-14
C118 4428 4541 4.46878e-15
C117 4429 4541 8.54023e-15
C116 4430 4541 1.11601e-14
C115 4431 4541 7.19482e-15
C114 4432 4541 7.37786e-15
C113 4433 4541 9.78565e-15
C112 4434 4541 1.57304e-14
C111 4435 4541 1.063e-14
C110 4436 4541 8.54023e-15
C109 4437 4541 1.11601e-14
C108 4438 4541 7.19482e-15
C107 4439 4541 4.46878e-15
C106 4440 4541 7.37786e-15
C105 4441 4541 9.78565e-15
C104 4442 4541 1.57304e-14
C103 4443 4541 1.063e-14
C102 4444 4541 3.45392e-14
C101 4445 4541 3.45392e-14
C100 4446 4541 3.45392e-14
C99 4447 4541 7.19482e-15
C98 4448 4541 4.46878e-15
C97 4449 4541 7.37786e-15
C96 4450 4541 9.78565e-15
C95 4451 4541 1.57304e-14
C94 4452 4541 4.78631e-14
C93 4453 4541 4.46878e-15
C92 4454 4541 7.19482e-15
C91 4455 4541 7.37786e-15
C90 4456 4541 9.78565e-15
C89 4457 4541 1.57304e-14
C88 4458 4541 6.59614e-14
C87 4459 4541 7.19482e-15
C86 4460 4541 4.46878e-15
C85 4461 4541 7.37786e-15
C84 4462 4541 9.78565e-15
C83 4463 4541 1.57304e-14
C82 4464 4541 6.89244e-14
C81 4465 4541 7.19482e-15
C80 4466 4541 4.46878e-15
C79 4467 4541 7.37786e-15
C78 4468 4541 9.78565e-15
C77 4469 4541 1.57304e-14
C76 4470 4541 7.93093e-14
C75 4471 4541 8.10579e-15
C74 4472 4541 8.10579e-15
C73 4473 4541 8.10579e-15
C72 4474 4541 8.10579e-15
C71 4475 4541 8.10579e-15
C70 4476 4541 8.18538e-13
C69 4477 4541 8.10579e-15
C68 4478 4541 1.59389e-11
C67 4479 4541 2.00607e-14
C66 4480 4541 1.84602e-14
C65 4481 4541 1.84602e-14
C64 4482 4541 2.00607e-14
C63 4483 4541 1.84602e-14
C62 4484 4541 2.00607e-14
C61 4485 4541 2.00607e-14
C60 4486 4541 1.84602e-14
C59 4487 4541 2.00607e-14
C58 4488 4541 1.84602e-14
C57 4489 4541 1.84602e-14
C56 4490 4541 2.00607e-14
C55 4491 4541 2.00607e-14
C54 4492 4541 1.84602e-14
C53 4493 4541 2.00607e-14
C52 4494 4541 1.84602e-14
C51 4495 4541 3.43699e-14
C50 4496 4541 2.1722e-14
C49 4497 4541 1.75135e-14
C48 4498 4541 1.91459e-14
C47 4499 4541 4.77843e-14
C46 4500 4541 3.43699e-14
C45 4501 4541 1.75135e-14
C44 4502 4541 2.1722e-14
C43 4503 4541 1.91459e-14
C42 4504 4541 4.77844e-14
C41 4505 4541 3.43699e-14
C40 4506 4541 1.75135e-14
C39 4507 4541 2.1722e-14
C38 4508 4541 1.91459e-14
C37 4509 4541 4.77843e-14
C36 4510 4541 3.43699e-14
C35 4511 4541 2.1722e-14
C34 4512 4541 1.75135e-14
C33 4513 4541 1.91459e-14
C32 4514 4541 4.77843e-14
C31 4515 4541 3.43699e-14
C30 4516 4541 2.1722e-14
C29 4517 4541 1.75135e-14
C28 4518 4541 1.91459e-14
C27 4519 4541 5.71705e-14
C26 4520 4541 3.43699e-14
C25 4521 4541 2.1722e-14
C24 4522 4541 1.75135e-14
C23 4523 4541 1.91459e-14
C22 4524 4541 5.71705e-14
C21 4525 4541 3.43699e-14
C20 4526 4541 1.75135e-14
C19 4527 4541 2.1722e-14
C18 4528 4541 1.91459e-14
C17 4529 4541 5.71705e-14
C16 4530 4541 3.43699e-14
C15 4531 4541 2.1722e-14
C14 4532 4541 1.75135e-14
C13 4533 4541 1.91459e-14
C12 4534 4541 5.71705e-14
C11 4535 4541 8.36649e-12
C10 4536 4541 1.77803e-13
C9 4537 4541 1.77803e-13
C8 4538 4541 1.77803e-13
C7 4539 4541 1.77803e-13
C6 4540 4541 1.53657e-11
C5 4541 4541 1.05845e-11
C4 4542 4541 1.87984e-13
C3 4543 4541 1.87984e-13
C2 4544 4541 1.87984e-13
C1 4545 4541 1.87984e-13
.ends amd2901

